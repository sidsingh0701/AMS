
module update_1 ( X, Y, Y_ramX, Y_ramY );
  input [15:0] X;
  input [15:0] Y;
  output [10:0] Y_ramX;
  output [10:0] Y_ramY;


  BUF_X4 U1 ( .A(X[4]), .Z(Y_ramX[0]) );
  BUF_X4 U2 ( .A(X[5]), .Z(Y_ramX[1]) );
  BUF_X4 U3 ( .A(X[6]), .Z(Y_ramX[2]) );
  BUF_X4 U4 ( .A(X[7]), .Z(Y_ramX[3]) );
  BUF_X4 U5 ( .A(X[8]), .Z(Y_ramX[4]) );
  BUF_X4 U6 ( .A(X[9]), .Z(Y_ramX[5]) );
  BUF_X4 U7 ( .A(X[10]), .Z(Y_ramX[6]) );
  BUF_X4 U8 ( .A(X[11]), .Z(Y_ramX[7]) );
  BUF_X4 U9 ( .A(X[12]), .Z(Y_ramX[8]) );
  BUF_X4 U10 ( .A(X[13]), .Z(Y_ramX[9]) );
  BUF_X4 U11 ( .A(X[14]), .Z(Y_ramX[10]) );
  BUF_X4 U12 ( .A(Y[8]), .Z(Y_ramY[4]) );
  BUF_X4 U13 ( .A(Y[9]), .Z(Y_ramY[5]) );
  BUF_X4 U14 ( .A(Y[10]), .Z(Y_ramY[6]) );
  BUF_X4 U15 ( .A(Y[11]), .Z(Y_ramY[7]) );
  BUF_X4 U16 ( .A(Y[12]), .Z(Y_ramY[8]) );
  BUF_X4 U17 ( .A(Y[13]), .Z(Y_ramY[9]) );
  BUF_X4 U18 ( .A(Y[14]), .Z(Y_ramY[10]) );
  BUF_X4 U19 ( .A(Y[4]), .Z(Y_ramY[0]) );
  BUF_X4 U20 ( .A(Y[5]), .Z(Y_ramY[1]) );
  BUF_X4 U21 ( .A(Y[6]), .Z(Y_ramY[2]) );
  BUF_X4 U22 ( .A(Y[7]), .Z(Y_ramY[3]) );
endmodule


module update_2 ( X, Y, RowX, RowY, Y_ramX, Y_ramY, Row_noX, Row_noY, clock, 
        EnableChange, FoundX, FoundY, FlagX, FlagY, DiagonalDoneX, 
        DiagonalDoneY, WireX, WireY );
  input [15:0] X;
  input [15:0] Y;
  input [255:0] RowX;
  input [255:0] RowY;
  input [10:0] Y_ramX;
  input [10:0] Y_ramY;
  output [10:0] Row_noX;
  output [10:0] Row_noY;
  input [1:0] FoundX;
  input [1:0] FoundY;
  input clock, EnableChange, FlagX, FlagY, DiagonalDoneX, DiagonalDoneY, WireX,
         WireY;
  wire   \U9/DATA16_0 , \U9/DATA16_1 , \U9/DATA16_2 , \U9/DATA16_3 ,
         \U9/DATA16_4 , \U9/DATA16_5 , \U9/DATA16_6 , \U9/DATA16_7 ,
         \U9/DATA16_8 , \U9/DATA16_9 , \U9/DATA16_10 , \U9/DATA15_0 ,
         \U9/DATA15_1 , \U9/DATA15_2 , \U9/DATA15_3 , \U9/DATA15_4 ,
         \U9/DATA15_5 , \U9/DATA15_6 , \U9/DATA15_7 , \U9/DATA15_8 ,
         \U9/DATA15_9 , \U9/DATA15_10 , \U9/DATA14_0 , \U9/DATA14_1 ,
         \U9/DATA14_2 , \U9/DATA14_3 , \U9/DATA14_4 , \U9/DATA14_5 ,
         \U9/DATA14_6 , \U9/DATA14_7 , \U9/DATA14_8 , \U9/DATA14_9 ,
         \U9/DATA14_10 , \U9/DATA13_0 , \U9/DATA13_1 , \U9/DATA13_2 ,
         \U9/DATA13_3 , \U9/DATA13_4 , \U9/DATA13_5 , \U9/DATA13_6 ,
         \U9/DATA13_7 , \U9/DATA13_8 , \U9/DATA13_9 , \U9/DATA13_10 ,
         \U9/DATA12_0 , \U9/DATA12_1 , \U9/DATA12_2 , \U9/DATA12_3 ,
         \U9/DATA12_4 , \U9/DATA12_5 , \U9/DATA12_6 , \U9/DATA12_7 ,
         \U9/DATA12_8 , \U9/DATA12_9 , \U9/DATA12_10 , \U9/DATA11_0 ,
         \U9/DATA11_1 , \U9/DATA11_2 , \U9/DATA11_3 , \U9/DATA11_4 ,
         \U9/DATA11_5 , \U9/DATA11_6 , \U9/DATA11_7 , \U9/DATA11_8 ,
         \U9/DATA11_9 , \U9/DATA11_10 , \U9/DATA10_0 , \U9/DATA10_1 ,
         \U9/DATA10_2 , \U9/DATA10_3 , \U9/DATA10_4 , \U9/DATA10_5 ,
         \U9/DATA10_6 , \U9/DATA10_7 , \U9/DATA10_8 , \U9/DATA10_9 ,
         \U9/DATA10_10 , \U9/DATA9_0 , \U9/DATA9_1 , \U9/DATA9_2 ,
         \U9/DATA9_3 , \U9/DATA9_4 , \U9/DATA9_5 , \U9/DATA9_6 , \U9/DATA9_7 ,
         \U9/DATA9_8 , \U9/DATA9_9 , \U9/DATA9_10 , \U9/DATA8_0 , \U9/DATA8_1 ,
         \U9/DATA8_2 , \U9/DATA8_3 , \U9/DATA8_4 , \U9/DATA8_5 , \U9/DATA8_6 ,
         \U9/DATA8_7 , \U9/DATA8_8 , \U9/DATA8_9 , \U9/DATA8_10 , \U9/DATA7_0 ,
         \U9/DATA7_1 , \U9/DATA7_2 , \U9/DATA7_3 , \U9/DATA7_4 , \U9/DATA7_5 ,
         \U9/DATA7_6 , \U9/DATA7_7 , \U9/DATA7_8 , \U9/DATA7_9 , \U9/DATA7_10 ,
         \U9/DATA6_0 , \U9/DATA6_1 , \U9/DATA6_2 , \U9/DATA6_3 , \U9/DATA6_4 ,
         \U9/DATA6_5 , \U9/DATA6_6 , \U9/DATA6_7 , \U9/DATA6_8 , \U9/DATA6_9 ,
         \U9/DATA6_10 , \U9/DATA5_0 , \U9/DATA5_1 , \U9/DATA5_2 , \U9/DATA5_3 ,
         \U9/DATA5_4 , \U9/DATA5_5 , \U9/DATA5_6 , \U9/DATA5_7 , \U9/DATA5_8 ,
         \U9/DATA5_9 , \U9/DATA5_10 , \U9/DATA4_0 , \U9/DATA4_1 , \U9/DATA4_2 ,
         \U9/DATA4_3 , \U9/DATA4_4 , \U9/DATA4_5 , \U9/DATA4_6 , \U9/DATA4_7 ,
         \U9/DATA4_8 , \U9/DATA4_9 , \U9/DATA4_10 , \U9/DATA3_0 , \U9/DATA3_1 ,
         \U9/DATA3_2 , \U9/DATA3_3 , \U9/DATA3_4 , \U9/DATA3_5 , \U9/DATA3_6 ,
         \U9/DATA3_7 , \U9/DATA3_8 , \U9/DATA3_9 , \U9/DATA3_10 , \U9/DATA2_0 ,
         \U9/DATA2_1 , \U9/DATA2_2 , \U9/DATA2_3 , \U9/DATA2_4 , \U9/DATA2_5 ,
         \U9/DATA2_6 , \U9/DATA2_7 , \U9/DATA2_8 , \U9/DATA2_9 , \U9/DATA2_10 ,
         \U9/DATA1_0 , \U9/DATA1_1 , \U9/DATA1_2 , \U9/DATA1_3 , \U9/DATA1_4 ,
         \U9/DATA1_5 , \U9/DATA1_6 , \U9/DATA1_7 , \U9/DATA1_8 , \U9/DATA1_9 ,
         \U9/DATA1_10 , \U8/DATA16_0 , \U8/DATA16_1 , \U8/DATA16_2 ,
         \U8/DATA16_3 , \U8/DATA16_4 , \U8/DATA16_5 , \U8/DATA16_6 ,
         \U8/DATA16_7 , \U8/DATA16_8 , \U8/DATA16_9 , \U8/DATA16_10 ,
         \U8/DATA15_0 , \U8/DATA15_1 , \U8/DATA15_2 , \U8/DATA15_3 ,
         \U8/DATA15_4 , \U8/DATA15_5 , \U8/DATA15_6 , \U8/DATA15_7 ,
         \U8/DATA15_8 , \U8/DATA15_9 , \U8/DATA15_10 , \U8/DATA14_0 ,
         \U8/DATA14_1 , \U8/DATA14_2 , \U8/DATA14_3 , \U8/DATA14_4 ,
         \U8/DATA14_5 , \U8/DATA14_6 , \U8/DATA14_7 , \U8/DATA14_8 ,
         \U8/DATA14_9 , \U8/DATA14_10 , \U8/DATA13_0 , \U8/DATA13_1 ,
         \U8/DATA13_2 , \U8/DATA13_3 , \U8/DATA13_4 , \U8/DATA13_5 ,
         \U8/DATA13_6 , \U8/DATA13_7 , \U8/DATA13_8 , \U8/DATA13_9 ,
         \U8/DATA13_10 , \U8/DATA12_0 , \U8/DATA12_1 , \U8/DATA12_2 ,
         \U8/DATA12_3 , \U8/DATA12_4 , \U8/DATA12_5 , \U8/DATA12_6 ,
         \U8/DATA12_7 , \U8/DATA12_8 , \U8/DATA12_9 , \U8/DATA12_10 ,
         \U8/DATA11_0 , \U8/DATA11_1 , \U8/DATA11_2 , \U8/DATA11_3 ,
         \U8/DATA11_4 , \U8/DATA11_5 , \U8/DATA11_6 , \U8/DATA11_7 ,
         \U8/DATA11_8 , \U8/DATA11_9 , \U8/DATA11_10 , \U8/DATA10_0 ,
         \U8/DATA10_1 , \U8/DATA10_2 , \U8/DATA10_3 , \U8/DATA10_4 ,
         \U8/DATA10_5 , \U8/DATA10_6 , \U8/DATA10_7 , \U8/DATA10_8 ,
         \U8/DATA10_9 , \U8/DATA10_10 , \U8/DATA9_0 , \U8/DATA9_1 ,
         \U8/DATA9_2 , \U8/DATA9_3 , \U8/DATA9_4 , \U8/DATA9_5 , \U8/DATA9_6 ,
         \U8/DATA9_7 , \U8/DATA9_8 , \U8/DATA9_9 , \U8/DATA9_10 , \U8/DATA8_0 ,
         \U8/DATA8_1 , \U8/DATA8_2 , \U8/DATA8_3 , \U8/DATA8_4 , \U8/DATA8_5 ,
         \U8/DATA8_6 , \U8/DATA8_7 , \U8/DATA8_8 , \U8/DATA8_9 , \U8/DATA8_10 ,
         \U8/DATA7_0 , \U8/DATA7_1 , \U8/DATA7_2 , \U8/DATA7_3 , \U8/DATA7_4 ,
         \U8/DATA7_5 , \U8/DATA7_6 , \U8/DATA7_7 , \U8/DATA7_8 , \U8/DATA7_9 ,
         \U8/DATA7_10 , \U8/DATA6_0 , \U8/DATA6_1 , \U8/DATA6_2 , \U8/DATA6_3 ,
         \U8/DATA6_4 , \U8/DATA6_5 , \U8/DATA6_6 , \U8/DATA6_7 , \U8/DATA6_8 ,
         \U8/DATA6_9 , \U8/DATA6_10 , \U8/DATA5_0 , \U8/DATA5_1 , \U8/DATA5_2 ,
         \U8/DATA5_3 , \U8/DATA5_4 , \U8/DATA5_5 , \U8/DATA5_6 , \U8/DATA5_7 ,
         \U8/DATA5_8 , \U8/DATA5_9 , \U8/DATA5_10 , \U8/DATA4_0 , \U8/DATA4_1 ,
         \U8/DATA4_2 , \U8/DATA4_3 , \U8/DATA4_4 , \U8/DATA4_5 , \U8/DATA4_6 ,
         \U8/DATA4_7 , \U8/DATA4_8 , \U8/DATA4_9 , \U8/DATA4_10 , \U8/DATA3_0 ,
         \U8/DATA3_1 , \U8/DATA3_2 , \U8/DATA3_3 , \U8/DATA3_4 , \U8/DATA3_5 ,
         \U8/DATA3_6 , \U8/DATA3_7 , \U8/DATA3_8 , \U8/DATA3_9 , \U8/DATA3_10 ,
         \U8/DATA2_0 , \U8/DATA2_1 , \U8/DATA2_2 , \U8/DATA2_3 , \U8/DATA2_4 ,
         \U8/DATA2_5 , \U8/DATA2_6 , \U8/DATA2_7 , \U8/DATA2_8 , \U8/DATA2_9 ,
         \U8/DATA2_10 , \U8/DATA1_0 , \U8/DATA1_1 , \U8/DATA1_2 , \U8/DATA1_3 ,
         \U8/DATA1_4 , \U8/DATA1_5 , \U8/DATA1_6 , \U8/DATA1_7 , \U8/DATA1_8 ,
         \U8/DATA1_9 , \U8/DATA1_10 , \U5/DATA1_1 , \U5/DATA1_2 , \U5/DATA1_3 ,
         \U5/DATA1_4 , \U5/DATA1_5 , \U5/DATA1_6 , \U5/DATA1_7 , \U5/DATA1_8 ,
         \U5/DATA1_9 , \U4/DATA1_1 , \U4/DATA1_2 , \U4/DATA1_3 , \U4/DATA1_4 ,
         \U4/DATA1_5 , \U4/DATA1_6 , \U4/DATA1_7 , \U4/DATA1_8 , \U4/DATA1_9 ,
         \add_93/carry[10] , \add_93/carry[9] , \add_93/carry[8] ,
         \add_93/carry[7] , \add_93/carry[6] , \add_93/carry[5] ,
         \add_93/carry[4] , \add_93/carry[3] , \add_93/carry[2] ,
         \add_93/A[0] , \add_93/A[1] , \add_93/A[2] , \add_93/A[3] ,
         \add_93/A[4] , \add_93/A[5] , \add_93/A[6] , \add_93/A[7] ,
         \add_93/A[8] , \add_93/A[9] , \add_93/A[10] , \add_87/carry[10] ,
         \add_87/carry[9] , \add_87/carry[8] , \add_87/carry[7] ,
         \add_87/carry[6] , \add_87/carry[5] , \add_87/carry[4] ,
         \add_87/carry[3] , \add_87/carry[2] , \add_87/A[0] , \add_87/A[1] ,
         \add_87/A[2] , \add_87/A[3] , \add_87/A[4] , \add_87/A[5] ,
         \add_87/A[6] , \add_87/A[7] , \add_87/A[8] , \add_87/A[9] ,
         \add_87/A[10] , n1, n12, n13, n24, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843;
  assign \U9/DATA16_0  = RowX[0];
  assign \U9/DATA16_1  = RowX[1];
  assign \U9/DATA16_2  = RowX[2];
  assign \U9/DATA16_3  = RowX[3];
  assign \U9/DATA16_4  = RowX[4];
  assign \U9/DATA16_5  = RowX[5];
  assign \U9/DATA16_6  = RowX[6];
  assign \U9/DATA16_7  = RowX[7];
  assign \U9/DATA16_8  = RowX[8];
  assign \U9/DATA16_9  = RowX[9];
  assign \U9/DATA16_10  = RowX[10];
  assign \U9/DATA15_0  = RowX[16];
  assign \U9/DATA15_1  = RowX[17];
  assign \U9/DATA15_2  = RowX[18];
  assign \U9/DATA15_3  = RowX[19];
  assign \U9/DATA15_4  = RowX[20];
  assign \U9/DATA15_5  = RowX[21];
  assign \U9/DATA15_6  = RowX[22];
  assign \U9/DATA15_7  = RowX[23];
  assign \U9/DATA15_8  = RowX[24];
  assign \U9/DATA15_9  = RowX[25];
  assign \U9/DATA15_10  = RowX[26];
  assign \U9/DATA14_0  = RowX[32];
  assign \U9/DATA14_1  = RowX[33];
  assign \U9/DATA14_2  = RowX[34];
  assign \U9/DATA14_3  = RowX[35];
  assign \U9/DATA14_4  = RowX[36];
  assign \U9/DATA14_5  = RowX[37];
  assign \U9/DATA14_6  = RowX[38];
  assign \U9/DATA14_7  = RowX[39];
  assign \U9/DATA14_8  = RowX[40];
  assign \U9/DATA14_9  = RowX[41];
  assign \U9/DATA14_10  = RowX[42];
  assign \U9/DATA13_0  = RowX[48];
  assign \U9/DATA13_1  = RowX[49];
  assign \U9/DATA13_2  = RowX[50];
  assign \U9/DATA13_3  = RowX[51];
  assign \U9/DATA13_4  = RowX[52];
  assign \U9/DATA13_5  = RowX[53];
  assign \U9/DATA13_6  = RowX[54];
  assign \U9/DATA13_7  = RowX[55];
  assign \U9/DATA13_8  = RowX[56];
  assign \U9/DATA13_9  = RowX[57];
  assign \U9/DATA13_10  = RowX[58];
  assign \U9/DATA12_0  = RowX[64];
  assign \U9/DATA12_1  = RowX[65];
  assign \U9/DATA12_2  = RowX[66];
  assign \U9/DATA12_3  = RowX[67];
  assign \U9/DATA12_4  = RowX[68];
  assign \U9/DATA12_5  = RowX[69];
  assign \U9/DATA12_6  = RowX[70];
  assign \U9/DATA12_7  = RowX[71];
  assign \U9/DATA12_8  = RowX[72];
  assign \U9/DATA12_9  = RowX[73];
  assign \U9/DATA12_10  = RowX[74];
  assign \U9/DATA11_0  = RowX[80];
  assign \U9/DATA11_1  = RowX[81];
  assign \U9/DATA11_2  = RowX[82];
  assign \U9/DATA11_3  = RowX[83];
  assign \U9/DATA11_4  = RowX[84];
  assign \U9/DATA11_5  = RowX[85];
  assign \U9/DATA11_6  = RowX[86];
  assign \U9/DATA11_7  = RowX[87];
  assign \U9/DATA11_8  = RowX[88];
  assign \U9/DATA11_9  = RowX[89];
  assign \U9/DATA11_10  = RowX[90];
  assign \U9/DATA10_0  = RowX[96];
  assign \U9/DATA10_1  = RowX[97];
  assign \U9/DATA10_2  = RowX[98];
  assign \U9/DATA10_3  = RowX[99];
  assign \U9/DATA10_4  = RowX[100];
  assign \U9/DATA10_5  = RowX[101];
  assign \U9/DATA10_6  = RowX[102];
  assign \U9/DATA10_7  = RowX[103];
  assign \U9/DATA10_8  = RowX[104];
  assign \U9/DATA10_9  = RowX[105];
  assign \U9/DATA10_10  = RowX[106];
  assign \U9/DATA9_0  = RowX[112];
  assign \U9/DATA9_1  = RowX[113];
  assign \U9/DATA9_2  = RowX[114];
  assign \U9/DATA9_3  = RowX[115];
  assign \U9/DATA9_4  = RowX[116];
  assign \U9/DATA9_5  = RowX[117];
  assign \U9/DATA9_6  = RowX[118];
  assign \U9/DATA9_7  = RowX[119];
  assign \U9/DATA9_8  = RowX[120];
  assign \U9/DATA9_9  = RowX[121];
  assign \U9/DATA9_10  = RowX[122];
  assign \U9/DATA8_0  = RowX[128];
  assign \U9/DATA8_1  = RowX[129];
  assign \U9/DATA8_2  = RowX[130];
  assign \U9/DATA8_3  = RowX[131];
  assign \U9/DATA8_4  = RowX[132];
  assign \U9/DATA8_5  = RowX[133];
  assign \U9/DATA8_6  = RowX[134];
  assign \U9/DATA8_7  = RowX[135];
  assign \U9/DATA8_8  = RowX[136];
  assign \U9/DATA8_9  = RowX[137];
  assign \U9/DATA8_10  = RowX[138];
  assign \U9/DATA7_0  = RowX[144];
  assign \U9/DATA7_1  = RowX[145];
  assign \U9/DATA7_2  = RowX[146];
  assign \U9/DATA7_3  = RowX[147];
  assign \U9/DATA7_4  = RowX[148];
  assign \U9/DATA7_5  = RowX[149];
  assign \U9/DATA7_6  = RowX[150];
  assign \U9/DATA7_7  = RowX[151];
  assign \U9/DATA7_8  = RowX[152];
  assign \U9/DATA7_9  = RowX[153];
  assign \U9/DATA7_10  = RowX[154];
  assign \U9/DATA6_0  = RowX[160];
  assign \U9/DATA6_1  = RowX[161];
  assign \U9/DATA6_2  = RowX[162];
  assign \U9/DATA6_3  = RowX[163];
  assign \U9/DATA6_4  = RowX[164];
  assign \U9/DATA6_5  = RowX[165];
  assign \U9/DATA6_6  = RowX[166];
  assign \U9/DATA6_7  = RowX[167];
  assign \U9/DATA6_8  = RowX[168];
  assign \U9/DATA6_9  = RowX[169];
  assign \U9/DATA6_10  = RowX[170];
  assign \U9/DATA5_0  = RowX[176];
  assign \U9/DATA5_1  = RowX[177];
  assign \U9/DATA5_2  = RowX[178];
  assign \U9/DATA5_3  = RowX[179];
  assign \U9/DATA5_4  = RowX[180];
  assign \U9/DATA5_5  = RowX[181];
  assign \U9/DATA5_6  = RowX[182];
  assign \U9/DATA5_7  = RowX[183];
  assign \U9/DATA5_8  = RowX[184];
  assign \U9/DATA5_9  = RowX[185];
  assign \U9/DATA5_10  = RowX[186];
  assign \U9/DATA4_0  = RowX[192];
  assign \U9/DATA4_1  = RowX[193];
  assign \U9/DATA4_2  = RowX[194];
  assign \U9/DATA4_3  = RowX[195];
  assign \U9/DATA4_4  = RowX[196];
  assign \U9/DATA4_5  = RowX[197];
  assign \U9/DATA4_6  = RowX[198];
  assign \U9/DATA4_7  = RowX[199];
  assign \U9/DATA4_8  = RowX[200];
  assign \U9/DATA4_9  = RowX[201];
  assign \U9/DATA4_10  = RowX[202];
  assign \U9/DATA3_0  = RowX[208];
  assign \U9/DATA3_1  = RowX[209];
  assign \U9/DATA3_2  = RowX[210];
  assign \U9/DATA3_3  = RowX[211];
  assign \U9/DATA3_4  = RowX[212];
  assign \U9/DATA3_5  = RowX[213];
  assign \U9/DATA3_6  = RowX[214];
  assign \U9/DATA3_7  = RowX[215];
  assign \U9/DATA3_8  = RowX[216];
  assign \U9/DATA3_9  = RowX[217];
  assign \U9/DATA3_10  = RowX[218];
  assign \U9/DATA2_0  = RowX[224];
  assign \U9/DATA2_1  = RowX[225];
  assign \U9/DATA2_2  = RowX[226];
  assign \U9/DATA2_3  = RowX[227];
  assign \U9/DATA2_4  = RowX[228];
  assign \U9/DATA2_5  = RowX[229];
  assign \U9/DATA2_6  = RowX[230];
  assign \U9/DATA2_7  = RowX[231];
  assign \U9/DATA2_8  = RowX[232];
  assign \U9/DATA2_9  = RowX[233];
  assign \U9/DATA2_10  = RowX[234];
  assign \U9/DATA1_0  = RowX[240];
  assign \U9/DATA1_1  = RowX[241];
  assign \U9/DATA1_2  = RowX[242];
  assign \U9/DATA1_3  = RowX[243];
  assign \U9/DATA1_4  = RowX[244];
  assign \U9/DATA1_5  = RowX[245];
  assign \U9/DATA1_6  = RowX[246];
  assign \U9/DATA1_7  = RowX[247];
  assign \U9/DATA1_8  = RowX[248];
  assign \U9/DATA1_9  = RowX[249];
  assign \U9/DATA1_10  = RowX[250];
  assign \U8/DATA16_0  = RowY[0];
  assign \U8/DATA16_1  = RowY[1];
  assign \U8/DATA16_2  = RowY[2];
  assign \U8/DATA16_3  = RowY[3];
  assign \U8/DATA16_4  = RowY[4];
  assign \U8/DATA16_5  = RowY[5];
  assign \U8/DATA16_6  = RowY[6];
  assign \U8/DATA16_7  = RowY[7];
  assign \U8/DATA16_8  = RowY[8];
  assign \U8/DATA16_9  = RowY[9];
  assign \U8/DATA16_10  = RowY[10];
  assign \U8/DATA15_0  = RowY[16];
  assign \U8/DATA15_1  = RowY[17];
  assign \U8/DATA15_2  = RowY[18];
  assign \U8/DATA15_3  = RowY[19];
  assign \U8/DATA15_4  = RowY[20];
  assign \U8/DATA15_5  = RowY[21];
  assign \U8/DATA15_6  = RowY[22];
  assign \U8/DATA15_7  = RowY[23];
  assign \U8/DATA15_8  = RowY[24];
  assign \U8/DATA15_9  = RowY[25];
  assign \U8/DATA15_10  = RowY[26];
  assign \U8/DATA14_0  = RowY[32];
  assign \U8/DATA14_1  = RowY[33];
  assign \U8/DATA14_2  = RowY[34];
  assign \U8/DATA14_3  = RowY[35];
  assign \U8/DATA14_4  = RowY[36];
  assign \U8/DATA14_5  = RowY[37];
  assign \U8/DATA14_6  = RowY[38];
  assign \U8/DATA14_7  = RowY[39];
  assign \U8/DATA14_8  = RowY[40];
  assign \U8/DATA14_9  = RowY[41];
  assign \U8/DATA14_10  = RowY[42];
  assign \U8/DATA13_0  = RowY[48];
  assign \U8/DATA13_1  = RowY[49];
  assign \U8/DATA13_2  = RowY[50];
  assign \U8/DATA13_3  = RowY[51];
  assign \U8/DATA13_4  = RowY[52];
  assign \U8/DATA13_5  = RowY[53];
  assign \U8/DATA13_6  = RowY[54];
  assign \U8/DATA13_7  = RowY[55];
  assign \U8/DATA13_8  = RowY[56];
  assign \U8/DATA13_9  = RowY[57];
  assign \U8/DATA13_10  = RowY[58];
  assign \U8/DATA12_0  = RowY[64];
  assign \U8/DATA12_1  = RowY[65];
  assign \U8/DATA12_2  = RowY[66];
  assign \U8/DATA12_3  = RowY[67];
  assign \U8/DATA12_4  = RowY[68];
  assign \U8/DATA12_5  = RowY[69];
  assign \U8/DATA12_6  = RowY[70];
  assign \U8/DATA12_7  = RowY[71];
  assign \U8/DATA12_8  = RowY[72];
  assign \U8/DATA12_9  = RowY[73];
  assign \U8/DATA12_10  = RowY[74];
  assign \U8/DATA11_0  = RowY[80];
  assign \U8/DATA11_1  = RowY[81];
  assign \U8/DATA11_2  = RowY[82];
  assign \U8/DATA11_3  = RowY[83];
  assign \U8/DATA11_4  = RowY[84];
  assign \U8/DATA11_5  = RowY[85];
  assign \U8/DATA11_6  = RowY[86];
  assign \U8/DATA11_7  = RowY[87];
  assign \U8/DATA11_8  = RowY[88];
  assign \U8/DATA11_9  = RowY[89];
  assign \U8/DATA11_10  = RowY[90];
  assign \U8/DATA10_0  = RowY[96];
  assign \U8/DATA10_1  = RowY[97];
  assign \U8/DATA10_2  = RowY[98];
  assign \U8/DATA10_3  = RowY[99];
  assign \U8/DATA10_4  = RowY[100];
  assign \U8/DATA10_5  = RowY[101];
  assign \U8/DATA10_6  = RowY[102];
  assign \U8/DATA10_7  = RowY[103];
  assign \U8/DATA10_8  = RowY[104];
  assign \U8/DATA10_9  = RowY[105];
  assign \U8/DATA10_10  = RowY[106];
  assign \U8/DATA9_0  = RowY[112];
  assign \U8/DATA9_1  = RowY[113];
  assign \U8/DATA9_2  = RowY[114];
  assign \U8/DATA9_3  = RowY[115];
  assign \U8/DATA9_4  = RowY[116];
  assign \U8/DATA9_5  = RowY[117];
  assign \U8/DATA9_6  = RowY[118];
  assign \U8/DATA9_7  = RowY[119];
  assign \U8/DATA9_8  = RowY[120];
  assign \U8/DATA9_9  = RowY[121];
  assign \U8/DATA9_10  = RowY[122];
  assign \U8/DATA8_0  = RowY[128];
  assign \U8/DATA8_1  = RowY[129];
  assign \U8/DATA8_2  = RowY[130];
  assign \U8/DATA8_3  = RowY[131];
  assign \U8/DATA8_4  = RowY[132];
  assign \U8/DATA8_5  = RowY[133];
  assign \U8/DATA8_6  = RowY[134];
  assign \U8/DATA8_7  = RowY[135];
  assign \U8/DATA8_8  = RowY[136];
  assign \U8/DATA8_9  = RowY[137];
  assign \U8/DATA8_10  = RowY[138];
  assign \U8/DATA7_0  = RowY[144];
  assign \U8/DATA7_1  = RowY[145];
  assign \U8/DATA7_2  = RowY[146];
  assign \U8/DATA7_3  = RowY[147];
  assign \U8/DATA7_4  = RowY[148];
  assign \U8/DATA7_5  = RowY[149];
  assign \U8/DATA7_6  = RowY[150];
  assign \U8/DATA7_7  = RowY[151];
  assign \U8/DATA7_8  = RowY[152];
  assign \U8/DATA7_9  = RowY[153];
  assign \U8/DATA7_10  = RowY[154];
  assign \U8/DATA6_0  = RowY[160];
  assign \U8/DATA6_1  = RowY[161];
  assign \U8/DATA6_2  = RowY[162];
  assign \U8/DATA6_3  = RowY[163];
  assign \U8/DATA6_4  = RowY[164];
  assign \U8/DATA6_5  = RowY[165];
  assign \U8/DATA6_6  = RowY[166];
  assign \U8/DATA6_7  = RowY[167];
  assign \U8/DATA6_8  = RowY[168];
  assign \U8/DATA6_9  = RowY[169];
  assign \U8/DATA6_10  = RowY[170];
  assign \U8/DATA5_0  = RowY[176];
  assign \U8/DATA5_1  = RowY[177];
  assign \U8/DATA5_2  = RowY[178];
  assign \U8/DATA5_3  = RowY[179];
  assign \U8/DATA5_4  = RowY[180];
  assign \U8/DATA5_5  = RowY[181];
  assign \U8/DATA5_6  = RowY[182];
  assign \U8/DATA5_7  = RowY[183];
  assign \U8/DATA5_8  = RowY[184];
  assign \U8/DATA5_9  = RowY[185];
  assign \U8/DATA5_10  = RowY[186];
  assign \U8/DATA4_0  = RowY[192];
  assign \U8/DATA4_1  = RowY[193];
  assign \U8/DATA4_2  = RowY[194];
  assign \U8/DATA4_3  = RowY[195];
  assign \U8/DATA4_4  = RowY[196];
  assign \U8/DATA4_5  = RowY[197];
  assign \U8/DATA4_6  = RowY[198];
  assign \U8/DATA4_7  = RowY[199];
  assign \U8/DATA4_8  = RowY[200];
  assign \U8/DATA4_9  = RowY[201];
  assign \U8/DATA4_10  = RowY[202];
  assign \U8/DATA3_0  = RowY[208];
  assign \U8/DATA3_1  = RowY[209];
  assign \U8/DATA3_2  = RowY[210];
  assign \U8/DATA3_3  = RowY[211];
  assign \U8/DATA3_4  = RowY[212];
  assign \U8/DATA3_5  = RowY[213];
  assign \U8/DATA3_6  = RowY[214];
  assign \U8/DATA3_7  = RowY[215];
  assign \U8/DATA3_8  = RowY[216];
  assign \U8/DATA3_9  = RowY[217];
  assign \U8/DATA3_10  = RowY[218];
  assign \U8/DATA2_0  = RowY[224];
  assign \U8/DATA2_1  = RowY[225];
  assign \U8/DATA2_2  = RowY[226];
  assign \U8/DATA2_3  = RowY[227];
  assign \U8/DATA2_4  = RowY[228];
  assign \U8/DATA2_5  = RowY[229];
  assign \U8/DATA2_6  = RowY[230];
  assign \U8/DATA2_7  = RowY[231];
  assign \U8/DATA2_8  = RowY[232];
  assign \U8/DATA2_9  = RowY[233];
  assign \U8/DATA2_10  = RowY[234];
  assign \U8/DATA1_0  = RowY[240];
  assign \U8/DATA1_1  = RowY[241];
  assign \U8/DATA1_2  = RowY[242];
  assign \U8/DATA1_3  = RowY[243];
  assign \U8/DATA1_4  = RowY[244];
  assign \U8/DATA1_5  = RowY[245];
  assign \U8/DATA1_6  = RowY[246];
  assign \U8/DATA1_7  = RowY[247];
  assign \U8/DATA1_8  = RowY[248];
  assign \U8/DATA1_9  = RowY[249];
  assign \U8/DATA1_10  = RowY[250];
  assign Row_noY[0] = \add_93/A[0] ;
  assign Row_noY[1] = \add_93/A[1] ;
  assign Row_noY[2] = \add_93/A[2] ;
  assign Row_noY[3] = \add_93/A[3] ;
  assign Row_noY[4] = \add_93/A[4] ;
  assign Row_noY[5] = \add_93/A[5] ;
  assign Row_noY[6] = \add_93/A[6] ;
  assign Row_noY[7] = \add_93/A[7] ;
  assign Row_noY[8] = \add_93/A[8] ;
  assign Row_noY[9] = \add_93/A[9] ;
  assign Row_noY[10] = \add_93/A[10] ;
  assign Row_noX[0] = \add_87/A[0] ;
  assign Row_noX[1] = \add_87/A[1] ;
  assign Row_noX[2] = \add_87/A[2] ;
  assign Row_noX[3] = \add_87/A[3] ;
  assign Row_noX[4] = \add_87/A[4] ;
  assign Row_noX[5] = \add_87/A[5] ;
  assign Row_noX[6] = \add_87/A[6] ;
  assign Row_noX[7] = \add_87/A[7] ;
  assign Row_noX[8] = \add_87/A[8] ;
  assign Row_noX[9] = \add_87/A[9] ;
  assign Row_noX[10] = \add_87/A[10] ;

  HA_X1 \add_87/U1_1_1  ( .A(\add_87/A[1] ), .B(\add_87/A[0] ), .CO(
        \add_87/carry[2] ), .S(\U5/DATA1_1 ) );
  HA_X1 \add_87/U1_1_2  ( .A(\add_87/A[2] ), .B(\add_87/carry[2] ), .CO(
        \add_87/carry[3] ), .S(\U5/DATA1_2 ) );
  HA_X1 \add_87/U1_1_3  ( .A(\add_87/A[3] ), .B(\add_87/carry[3] ), .CO(
        \add_87/carry[4] ), .S(\U5/DATA1_3 ) );
  HA_X1 \add_87/U1_1_4  ( .A(\add_87/A[4] ), .B(\add_87/carry[4] ), .CO(
        \add_87/carry[5] ), .S(\U5/DATA1_4 ) );
  HA_X1 \add_87/U1_1_5  ( .A(\add_87/A[5] ), .B(\add_87/carry[5] ), .CO(
        \add_87/carry[6] ), .S(\U5/DATA1_5 ) );
  HA_X1 \add_87/U1_1_6  ( .A(\add_87/A[6] ), .B(\add_87/carry[6] ), .CO(
        \add_87/carry[7] ), .S(\U5/DATA1_6 ) );
  HA_X1 \add_87/U1_1_7  ( .A(\add_87/A[7] ), .B(\add_87/carry[7] ), .CO(
        \add_87/carry[8] ), .S(\U5/DATA1_7 ) );
  HA_X1 \add_87/U1_1_8  ( .A(\add_87/A[8] ), .B(\add_87/carry[8] ), .CO(
        \add_87/carry[9] ), .S(\U5/DATA1_8 ) );
  HA_X1 \add_87/U1_1_9  ( .A(\add_87/A[9] ), .B(\add_87/carry[9] ), .CO(
        \add_87/carry[10] ), .S(\U5/DATA1_9 ) );
  HA_X1 \add_93/U1_1_1  ( .A(\add_93/A[1] ), .B(\add_93/A[0] ), .CO(
        \add_93/carry[2] ), .S(\U4/DATA1_1 ) );
  HA_X1 \add_93/U1_1_2  ( .A(\add_93/A[2] ), .B(\add_93/carry[2] ), .CO(
        \add_93/carry[3] ), .S(\U4/DATA1_2 ) );
  HA_X1 \add_93/U1_1_3  ( .A(\add_93/A[3] ), .B(\add_93/carry[3] ), .CO(
        \add_93/carry[4] ), .S(\U4/DATA1_3 ) );
  HA_X1 \add_93/U1_1_4  ( .A(\add_93/A[4] ), .B(\add_93/carry[4] ), .CO(
        \add_93/carry[5] ), .S(\U4/DATA1_4 ) );
  HA_X1 \add_93/U1_1_5  ( .A(\add_93/A[5] ), .B(\add_93/carry[5] ), .CO(
        \add_93/carry[6] ), .S(\U4/DATA1_5 ) );
  HA_X1 \add_93/U1_1_6  ( .A(\add_93/A[6] ), .B(\add_93/carry[6] ), .CO(
        \add_93/carry[7] ), .S(\U4/DATA1_6 ) );
  HA_X1 \add_93/U1_1_7  ( .A(\add_93/A[7] ), .B(\add_93/carry[7] ), .CO(
        \add_93/carry[8] ), .S(\U4/DATA1_7 ) );
  HA_X1 \add_93/U1_1_8  ( .A(\add_93/A[8] ), .B(\add_93/carry[8] ), .CO(
        \add_93/carry[9] ), .S(\U4/DATA1_8 ) );
  HA_X1 \add_93/U1_1_9  ( .A(\add_93/A[9] ), .B(\add_93/carry[9] ), .CO(
        \add_93/carry[10] ), .S(\U4/DATA1_9 ) );
  DFF_X1 \Row_noX_reg[0]  ( .D(n365), .CK(clock), .Q(\add_87/A[0] ), .QN(n12)
         );
  DFF_X1 \Row_noX_reg[1]  ( .D(n830), .CK(clock), .Q(\add_87/A[1] ) );
  DFF_X1 \Row_noX_reg[2]  ( .D(n829), .CK(clock), .Q(\add_87/A[2] ) );
  DFF_X1 \Row_noX_reg[3]  ( .D(n828), .CK(clock), .Q(\add_87/A[3] ) );
  DFF_X1 \Row_noX_reg[4]  ( .D(n827), .CK(clock), .Q(\add_87/A[4] ) );
  DFF_X1 \Row_noX_reg[5]  ( .D(n826), .CK(clock), .Q(\add_87/A[5] ) );
  DFF_X1 \Row_noX_reg[6]  ( .D(n825), .CK(clock), .Q(\add_87/A[6] ) );
  DFF_X1 \Row_noX_reg[7]  ( .D(n824), .CK(clock), .Q(\add_87/A[7] ) );
  DFF_X1 \Row_noX_reg[8]  ( .D(n823), .CK(clock), .Q(\add_87/A[8] ) );
  DFF_X1 \Row_noX_reg[9]  ( .D(n822), .CK(clock), .Q(\add_87/A[9] ) );
  DFF_X1 \Row_noY_reg[0]  ( .D(n363), .CK(clock), .Q(\add_93/A[0] ), .QN(n24)
         );
  DFF_X1 \Row_noY_reg[1]  ( .D(n817), .CK(clock), .Q(\add_93/A[1] ) );
  DFF_X1 \Row_noY_reg[2]  ( .D(n816), .CK(clock), .Q(\add_93/A[2] ) );
  DFF_X1 \Row_noY_reg[3]  ( .D(n815), .CK(clock), .Q(\add_93/A[3] ) );
  DFF_X1 \Row_noY_reg[4]  ( .D(n814), .CK(clock), .Q(\add_93/A[4] ) );
  DFF_X1 \Row_noY_reg[5]  ( .D(n813), .CK(clock), .Q(\add_93/A[5] ) );
  DFF_X1 \Row_noY_reg[6]  ( .D(n812), .CK(clock), .Q(\add_93/A[6] ) );
  DFF_X1 \Row_noY_reg[7]  ( .D(n811), .CK(clock), .Q(\add_93/A[7] ) );
  DFF_X1 \Row_noY_reg[8]  ( .D(n810), .CK(clock), .Q(\add_93/A[8] ) );
  DFF_X1 \Row_noY_reg[9]  ( .D(n809), .CK(clock), .Q(\add_93/A[9] ) );
  NAND4_X2 U5 ( .A1(n45), .A2(n46), .A3(n47), .A4(n48), .ZN(n43) );
  NAND4_X2 U10 ( .A1(n57), .A2(n58), .A3(n59), .A4(n60), .ZN(n42) );
  NAND3_X2 U15 ( .A1(n819), .A2(n13), .A3(\add_93/carry[10] ), .ZN(n40) );
  AOI221_X2 U17 ( .B1(\add_93/A[9] ), .B2(n820), .C1(\U4/DATA1_9 ), .C2(n819), 
        .A(n73), .ZN(n72) );
  AND4_X2 U19 ( .A1(n76), .A2(n77), .A3(n78), .A4(n79), .ZN(n75) );
  AND4_X2 U24 ( .A1(n80), .A2(n81), .A3(n82), .A4(n83), .ZN(n74) );
  AOI221_X2 U29 ( .B1(\add_93/A[8] ), .B2(n820), .C1(\U4/DATA1_8 ), .C2(n819), 
        .A(n85), .ZN(n84) );
  AND4_X2 U31 ( .A1(n88), .A2(n89), .A3(n90), .A4(n91), .ZN(n87) );
  AND4_X2 U36 ( .A1(n92), .A2(n93), .A3(n94), .A4(n95), .ZN(n86) );
  AOI221_X2 U41 ( .B1(\add_93/A[7] ), .B2(n820), .C1(\U4/DATA1_7 ), .C2(n819), 
        .A(n97), .ZN(n96) );
  AND4_X2 U43 ( .A1(n100), .A2(n101), .A3(n102), .A4(n103), .ZN(n99) );
  AND4_X2 U48 ( .A1(n104), .A2(n105), .A3(n106), .A4(n107), .ZN(n98) );
  AOI221_X2 U53 ( .B1(\add_93/A[6] ), .B2(n820), .C1(\U4/DATA1_6 ), .C2(n819), 
        .A(n109), .ZN(n108) );
  AND4_X2 U55 ( .A1(n112), .A2(n113), .A3(n114), .A4(n115), .ZN(n111) );
  AND4_X2 U60 ( .A1(n116), .A2(n117), .A3(n118), .A4(n119), .ZN(n110) );
  AOI221_X2 U65 ( .B1(\add_93/A[5] ), .B2(n820), .C1(\U4/DATA1_5 ), .C2(n819), 
        .A(n121), .ZN(n120) );
  AND4_X2 U67 ( .A1(n124), .A2(n125), .A3(n126), .A4(n127), .ZN(n123) );
  AND4_X2 U72 ( .A1(n128), .A2(n129), .A3(n130), .A4(n131), .ZN(n122) );
  AOI221_X2 U77 ( .B1(\add_93/A[4] ), .B2(n820), .C1(\U4/DATA1_4 ), .C2(n819), 
        .A(n133), .ZN(n132) );
  AND4_X2 U79 ( .A1(n136), .A2(n137), .A3(n138), .A4(n139), .ZN(n135) );
  AND4_X2 U84 ( .A1(n140), .A2(n141), .A3(n142), .A4(n143), .ZN(n134) );
  AOI221_X2 U89 ( .B1(\add_93/A[3] ), .B2(n820), .C1(\U4/DATA1_3 ), .C2(n819), 
        .A(n145), .ZN(n144) );
  AND4_X2 U91 ( .A1(n148), .A2(n149), .A3(n150), .A4(n151), .ZN(n147) );
  AND4_X2 U96 ( .A1(n152), .A2(n153), .A3(n154), .A4(n155), .ZN(n146) );
  AOI221_X2 U101 ( .B1(\add_93/A[2] ), .B2(n820), .C1(\U4/DATA1_2 ), .C2(n819), 
        .A(n157), .ZN(n156) );
  AND4_X2 U103 ( .A1(n160), .A2(n161), .A3(n162), .A4(n163), .ZN(n159) );
  AND4_X2 U108 ( .A1(n164), .A2(n165), .A3(n166), .A4(n167), .ZN(n158) );
  AOI221_X2 U113 ( .B1(\add_93/A[1] ), .B2(n820), .C1(\U4/DATA1_1 ), .C2(n819), 
        .A(n169), .ZN(n168) );
  AND4_X2 U115 ( .A1(n172), .A2(n173), .A3(n174), .A4(n175), .ZN(n171) );
  AND4_X2 U120 ( .A1(n176), .A2(n177), .A3(n178), .A4(n179), .ZN(n170) );
  OAI221_X2 U125 ( .B1(\add_93/A[0] ), .B2(n70), .C1(n71), .C2(n24), .A(n180), 
        .ZN(n363) );
  NOR2_X2 U127 ( .A1(n819), .A2(n820), .ZN(n44) );
  NAND4_X2 U128 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(n182) );
  NOR2_X2 U133 ( .A1(Y[3]), .A2(Y[0]), .ZN(n187) );
  NOR2_X2 U134 ( .A1(n843), .A2(Y[3]), .ZN(n189) );
  NAND4_X2 U135 ( .A1(n193), .A2(n194), .A3(n195), .A4(n196), .ZN(n181) );
  NOR2_X2 U139 ( .A1(n842), .A2(Y[2]), .ZN(n191) );
  NOR2_X2 U141 ( .A1(n841), .A2(Y[0]), .ZN(n197) );
  NOR2_X2 U142 ( .A1(n841), .A2(n843), .ZN(n198) );
  NOR2_X2 U143 ( .A1(Y[2]), .A2(Y[1]), .ZN(n192) );
  NAND2_X2 U144 ( .A1(n70), .A2(n199), .ZN(n71) );
  NAND2_X2 U145 ( .A1(FlagY), .A2(n836), .ZN(n199) );
  NOR2_X2 U147 ( .A1(FoundY[1]), .A2(n836), .ZN(n200) );
  OAI221_X2 U148 ( .B1(n837), .B2(n201), .C1(n202), .C2(n1), .A(n203), .ZN(
        n364) );
  NAND4_X2 U150 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(n205) );
  NAND4_X2 U155 ( .A1(n219), .A2(n220), .A3(n221), .A4(n222), .ZN(n204) );
  NAND2_X2 U161 ( .A1(n832), .A2(n1), .ZN(n201) );
  AOI221_X2 U162 ( .B1(\add_87/A[9] ), .B2(n833), .C1(\U5/DATA1_9 ), .C2(n832), 
        .A(n232), .ZN(n231) );
  AND4_X2 U164 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(n234) );
  AND4_X2 U169 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(n233) );
  AOI221_X2 U174 ( .B1(\add_87/A[8] ), .B2(n833), .C1(\U5/DATA1_8 ), .C2(n832), 
        .A(n244), .ZN(n243) );
  AND4_X2 U176 ( .A1(n247), .A2(n248), .A3(n249), .A4(n250), .ZN(n246) );
  AND4_X2 U181 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(n245) );
  AOI221_X2 U186 ( .B1(\add_87/A[7] ), .B2(n833), .C1(\U5/DATA1_7 ), .C2(n832), 
        .A(n256), .ZN(n255) );
  AND4_X2 U188 ( .A1(n259), .A2(n260), .A3(n261), .A4(n262), .ZN(n258) );
  AND4_X2 U193 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(n257) );
  AOI221_X2 U198 ( .B1(\add_87/A[6] ), .B2(n833), .C1(\U5/DATA1_6 ), .C2(n832), 
        .A(n268), .ZN(n267) );
  AND4_X2 U200 ( .A1(n271), .A2(n272), .A3(n273), .A4(n274), .ZN(n270) );
  AND4_X2 U205 ( .A1(n275), .A2(n276), .A3(n277), .A4(n278), .ZN(n269) );
  AOI221_X2 U210 ( .B1(\add_87/A[5] ), .B2(n833), .C1(\U5/DATA1_5 ), .C2(n832), 
        .A(n280), .ZN(n279) );
  AND4_X2 U212 ( .A1(n283), .A2(n284), .A3(n285), .A4(n286), .ZN(n282) );
  AND4_X2 U217 ( .A1(n287), .A2(n288), .A3(n289), .A4(n290), .ZN(n281) );
  AOI221_X2 U222 ( .B1(\add_87/A[4] ), .B2(n833), .C1(\U5/DATA1_4 ), .C2(n832), 
        .A(n292), .ZN(n291) );
  AND4_X2 U224 ( .A1(n295), .A2(n296), .A3(n297), .A4(n298), .ZN(n294) );
  AND4_X2 U229 ( .A1(n299), .A2(n300), .A3(n301), .A4(n302), .ZN(n293) );
  AOI221_X2 U234 ( .B1(\add_87/A[3] ), .B2(n833), .C1(\U5/DATA1_3 ), .C2(n832), 
        .A(n304), .ZN(n303) );
  AND4_X2 U236 ( .A1(n307), .A2(n308), .A3(n309), .A4(n310), .ZN(n306) );
  AND4_X2 U241 ( .A1(n311), .A2(n312), .A3(n313), .A4(n314), .ZN(n305) );
  AOI221_X2 U246 ( .B1(\add_87/A[2] ), .B2(n833), .C1(\U5/DATA1_2 ), .C2(n832), 
        .A(n316), .ZN(n315) );
  AND4_X2 U248 ( .A1(n319), .A2(n320), .A3(n321), .A4(n322), .ZN(n318) );
  AND4_X2 U253 ( .A1(n323), .A2(n324), .A3(n325), .A4(n326), .ZN(n317) );
  AOI221_X2 U258 ( .B1(\add_87/A[1] ), .B2(n833), .C1(\U5/DATA1_1 ), .C2(n832), 
        .A(n328), .ZN(n327) );
  AND4_X2 U260 ( .A1(n331), .A2(n332), .A3(n333), .A4(n334), .ZN(n330) );
  AND4_X2 U265 ( .A1(n335), .A2(n336), .A3(n337), .A4(n338), .ZN(n329) );
  OAI221_X2 U270 ( .B1(\add_87/A[0] ), .B2(n339), .C1(n340), .C2(n12), .A(n341), .ZN(n365) );
  NOR2_X2 U272 ( .A1(n833), .A2(n832), .ZN(n206) );
  NAND4_X2 U273 ( .A1(n344), .A2(n345), .A3(n346), .A4(n347), .ZN(n343) );
  NOR2_X2 U278 ( .A1(X[3]), .A2(X[0]), .ZN(n348) );
  NOR2_X2 U279 ( .A1(n840), .A2(X[3]), .ZN(n350) );
  NAND4_X2 U280 ( .A1(n354), .A2(n355), .A3(n356), .A4(n357), .ZN(n342) );
  NOR2_X2 U284 ( .A1(n839), .A2(X[2]), .ZN(n352) );
  NOR2_X2 U286 ( .A1(n838), .A2(X[0]), .ZN(n358) );
  NOR2_X2 U287 ( .A1(n838), .A2(n840), .ZN(n359) );
  NOR2_X2 U288 ( .A1(X[2]), .A2(X[1]), .ZN(n353) );
  NAND2_X2 U289 ( .A1(n339), .A2(n360), .ZN(n340) );
  NAND2_X2 U290 ( .A1(FlagX), .A2(n835), .ZN(n360) );
  NOR2_X2 U292 ( .A1(FoundX[1]), .A2(n834), .ZN(n361) );
  AND2_X1 U338 ( .A1(Y[2]), .A2(Y[1]), .ZN(n188) );
  AND2_X1 U341 ( .A1(Y[2]), .A2(n842), .ZN(n190) );
  AND2_X1 U356 ( .A1(X[2]), .A2(X[1]), .ZN(n349) );
  AND2_X1 U359 ( .A1(X[2]), .A2(n839), .ZN(n351) );
  DFF_X2 \Row_noX_reg[10]  ( .D(n364), .CK(clock), .Q(\add_87/A[10] ), .QN(n1)
         );
  DFF_X2 \Row_noY_reg[10]  ( .D(n362), .CK(clock), .Q(\add_93/A[10] ), .QN(n13) );
  AOI22_X2 U3 ( .A1(\U8/DATA10_10 ), .A2(n67), .B1(\U8/DATA9_10 ), .B2(n68), 
        .ZN(n57) );
  AOI22_X2 U4 ( .A1(\U8/DATA12_10 ), .A2(n65), .B1(\U8/DATA11_10 ), .B2(n66), 
        .ZN(n58) );
  AOI22_X2 U6 ( .A1(\U8/DATA16_10 ), .A2(n61), .B1(\U8/DATA15_10 ), .B2(n62), 
        .ZN(n60) );
  AOI22_X2 U7 ( .A1(\U9/DATA10_10 ), .A2(n229), .B1(\U9/DATA9_10 ), .B2(n230), 
        .ZN(n219) );
  AOI22_X2 U8 ( .A1(\U9/DATA12_10 ), .A2(n227), .B1(\U9/DATA11_10 ), .B2(n228), 
        .ZN(n220) );
  AOI22_X2 U9 ( .A1(\U9/DATA16_10 ), .A2(n223), .B1(\U9/DATA15_10 ), .B2(n224), 
        .ZN(n222) );
  AOI22_X2 U11 ( .A1(\U9/DATA10_0 ), .A2(n229), .B1(\U9/DATA9_0 ), .B2(n230), 
        .ZN(n354) );
  AOI22_X2 U12 ( .A1(\U8/DATA2_10 ), .A2(n55), .B1(\U8/DATA1_10 ), .B2(n56), 
        .ZN(n45) );
  AOI22_X2 U13 ( .A1(\U8/DATA4_10 ), .A2(n53), .B1(\U8/DATA3_10 ), .B2(n54), 
        .ZN(n46) );
  AOI22_X2 U14 ( .A1(\U8/DATA8_10 ), .A2(n49), .B1(\U8/DATA7_10 ), .B2(n50), 
        .ZN(n48) );
  AOI22_X2 U16 ( .A1(\U9/DATA2_10 ), .A2(n217), .B1(\U9/DATA1_10 ), .B2(n218), 
        .ZN(n207) );
  AOI22_X2 U18 ( .A1(\U9/DATA4_10 ), .A2(n215), .B1(\U9/DATA3_10 ), .B2(n216), 
        .ZN(n208) );
  AOI22_X2 U20 ( .A1(\U9/DATA8_10 ), .A2(n211), .B1(\U9/DATA7_10 ), .B2(n212), 
        .ZN(n210) );
  AOI22_X2 U21 ( .A1(\U9/DATA12_0 ), .A2(n227), .B1(\U9/DATA11_0 ), .B2(n228), 
        .ZN(n355) );
  AOI22_X2 U22 ( .A1(\U9/DATA12_9 ), .A2(n227), .B1(\U9/DATA11_9 ), .B2(n228), 
        .ZN(n236) );
  AOI22_X2 U23 ( .A1(\U9/DATA12_8 ), .A2(n227), .B1(\U9/DATA11_8 ), .B2(n228), 
        .ZN(n248) );
  AOI22_X2 U25 ( .A1(\U9/DATA12_7 ), .A2(n227), .B1(\U9/DATA11_7 ), .B2(n228), 
        .ZN(n260) );
  AOI22_X2 U26 ( .A1(\U9/DATA12_6 ), .A2(n227), .B1(\U9/DATA11_6 ), .B2(n228), 
        .ZN(n272) );
  AOI22_X2 U27 ( .A1(\U9/DATA12_5 ), .A2(n227), .B1(\U9/DATA11_5 ), .B2(n228), 
        .ZN(n284) );
  AOI22_X2 U28 ( .A1(\U9/DATA12_4 ), .A2(n227), .B1(\U9/DATA11_4 ), .B2(n228), 
        .ZN(n296) );
  AOI22_X2 U30 ( .A1(\U9/DATA12_3 ), .A2(n227), .B1(\U9/DATA11_3 ), .B2(n228), 
        .ZN(n308) );
  AOI22_X2 U32 ( .A1(\U9/DATA12_2 ), .A2(n227), .B1(\U9/DATA11_2 ), .B2(n228), 
        .ZN(n320) );
  AOI22_X2 U33 ( .A1(\U9/DATA12_1 ), .A2(n227), .B1(\U9/DATA11_1 ), .B2(n228), 
        .ZN(n332) );
  AOI22_X2 U34 ( .A1(\U9/DATA10_9 ), .A2(n229), .B1(\U9/DATA9_9 ), .B2(n230), 
        .ZN(n235) );
  AOI22_X2 U35 ( .A1(\U9/DATA10_8 ), .A2(n229), .B1(\U9/DATA9_8 ), .B2(n230), 
        .ZN(n247) );
  AOI22_X2 U37 ( .A1(\U9/DATA10_7 ), .A2(n229), .B1(\U9/DATA9_7 ), .B2(n230), 
        .ZN(n259) );
  AOI22_X2 U38 ( .A1(\U9/DATA10_6 ), .A2(n229), .B1(\U9/DATA9_6 ), .B2(n230), 
        .ZN(n271) );
  AOI22_X2 U39 ( .A1(\U9/DATA10_5 ), .A2(n229), .B1(\U9/DATA9_5 ), .B2(n230), 
        .ZN(n283) );
  AOI22_X2 U40 ( .A1(\U9/DATA10_4 ), .A2(n229), .B1(\U9/DATA9_4 ), .B2(n230), 
        .ZN(n295) );
  AOI22_X2 U42 ( .A1(\U9/DATA10_3 ), .A2(n229), .B1(\U9/DATA9_3 ), .B2(n230), 
        .ZN(n307) );
  AOI22_X2 U44 ( .A1(\U9/DATA10_2 ), .A2(n229), .B1(\U9/DATA9_2 ), .B2(n230), 
        .ZN(n319) );
  AOI22_X2 U45 ( .A1(\U9/DATA10_1 ), .A2(n229), .B1(\U9/DATA9_1 ), .B2(n230), 
        .ZN(n331) );
  OAI21_X2 U46 ( .B1(n70), .B2(\add_93/carry[10] ), .A(n71), .ZN(n69) );
  AOI22_X2 U47 ( .A1(\U8/DATA8_9 ), .A2(n49), .B1(\U8/DATA7_9 ), .B2(n50), 
        .ZN(n83) );
  AOI22_X2 U49 ( .A1(\U8/DATA2_9 ), .A2(n55), .B1(\U8/DATA1_9 ), .B2(n56), 
        .ZN(n80) );
  AOI22_X2 U50 ( .A1(\U8/DATA4_9 ), .A2(n53), .B1(\U8/DATA3_9 ), .B2(n54), 
        .ZN(n81) );
  AOI22_X2 U51 ( .A1(\U8/DATA8_8 ), .A2(n49), .B1(\U8/DATA7_8 ), .B2(n50), 
        .ZN(n95) );
  AOI22_X2 U52 ( .A1(\U8/DATA2_8 ), .A2(n55), .B1(\U8/DATA1_8 ), .B2(n56), 
        .ZN(n92) );
  AOI22_X2 U54 ( .A1(\U8/DATA4_8 ), .A2(n53), .B1(\U8/DATA3_8 ), .B2(n54), 
        .ZN(n93) );
  AOI22_X2 U56 ( .A1(\U8/DATA8_7 ), .A2(n49), .B1(\U8/DATA7_7 ), .B2(n50), 
        .ZN(n107) );
  AOI22_X2 U57 ( .A1(\U8/DATA2_7 ), .A2(n55), .B1(\U8/DATA1_7 ), .B2(n56), 
        .ZN(n104) );
  AOI22_X2 U58 ( .A1(\U8/DATA4_7 ), .A2(n53), .B1(\U8/DATA3_7 ), .B2(n54), 
        .ZN(n105) );
  AOI22_X2 U59 ( .A1(\U8/DATA8_6 ), .A2(n49), .B1(\U8/DATA7_6 ), .B2(n50), 
        .ZN(n119) );
  AOI22_X2 U61 ( .A1(\U8/DATA2_6 ), .A2(n55), .B1(\U8/DATA1_6 ), .B2(n56), 
        .ZN(n116) );
  AOI22_X2 U62 ( .A1(\U8/DATA4_6 ), .A2(n53), .B1(\U8/DATA3_6 ), .B2(n54), 
        .ZN(n117) );
  AOI22_X2 U63 ( .A1(\U8/DATA8_5 ), .A2(n49), .B1(\U8/DATA7_5 ), .B2(n50), 
        .ZN(n131) );
  AOI22_X2 U64 ( .A1(\U8/DATA2_5 ), .A2(n55), .B1(\U8/DATA1_5 ), .B2(n56), 
        .ZN(n128) );
  AOI22_X2 U66 ( .A1(\U8/DATA4_5 ), .A2(n53), .B1(\U8/DATA3_5 ), .B2(n54), 
        .ZN(n129) );
  AOI22_X2 U68 ( .A1(\U8/DATA8_4 ), .A2(n49), .B1(\U8/DATA7_4 ), .B2(n50), 
        .ZN(n143) );
  AOI22_X2 U69 ( .A1(\U8/DATA2_4 ), .A2(n55), .B1(\U8/DATA1_4 ), .B2(n56), 
        .ZN(n140) );
  AOI22_X2 U70 ( .A1(\U8/DATA4_4 ), .A2(n53), .B1(\U8/DATA3_4 ), .B2(n54), 
        .ZN(n141) );
  AOI22_X2 U71 ( .A1(\U8/DATA8_3 ), .A2(n49), .B1(\U8/DATA7_3 ), .B2(n50), 
        .ZN(n155) );
  AOI22_X2 U73 ( .A1(\U8/DATA2_3 ), .A2(n55), .B1(\U8/DATA1_3 ), .B2(n56), 
        .ZN(n152) );
  AOI22_X2 U74 ( .A1(\U8/DATA4_3 ), .A2(n53), .B1(\U8/DATA3_3 ), .B2(n54), 
        .ZN(n153) );
  AOI22_X2 U75 ( .A1(\U8/DATA8_2 ), .A2(n49), .B1(\U8/DATA7_2 ), .B2(n50), 
        .ZN(n167) );
  AOI22_X2 U76 ( .A1(\U8/DATA2_2 ), .A2(n55), .B1(\U8/DATA1_2 ), .B2(n56), 
        .ZN(n164) );
  AOI22_X2 U78 ( .A1(\U8/DATA4_2 ), .A2(n53), .B1(\U8/DATA3_2 ), .B2(n54), 
        .ZN(n165) );
  AOI22_X2 U80 ( .A1(\U8/DATA8_1 ), .A2(n49), .B1(\U8/DATA7_1 ), .B2(n50), 
        .ZN(n179) );
  AOI22_X2 U81 ( .A1(\U8/DATA2_1 ), .A2(n55), .B1(\U8/DATA1_1 ), .B2(n56), 
        .ZN(n176) );
  AOI22_X2 U82 ( .A1(\U8/DATA4_1 ), .A2(n53), .B1(\U8/DATA3_1 ), .B2(n54), 
        .ZN(n177) );
  AOI22_X2 U83 ( .A1(\U9/DATA8_9 ), .A2(n211), .B1(\U9/DATA7_9 ), .B2(n212), 
        .ZN(n242) );
  AOI22_X2 U85 ( .A1(\U9/DATA2_9 ), .A2(n217), .B1(\U9/DATA1_9 ), .B2(n218), 
        .ZN(n239) );
  AOI22_X2 U86 ( .A1(\U9/DATA4_9 ), .A2(n215), .B1(\U9/DATA3_9 ), .B2(n216), 
        .ZN(n240) );
  AOI22_X2 U87 ( .A1(\U9/DATA8_8 ), .A2(n211), .B1(\U9/DATA7_8 ), .B2(n212), 
        .ZN(n254) );
  AOI22_X2 U88 ( .A1(\U9/DATA2_8 ), .A2(n217), .B1(\U9/DATA1_8 ), .B2(n218), 
        .ZN(n251) );
  AOI22_X2 U90 ( .A1(\U9/DATA4_8 ), .A2(n215), .B1(\U9/DATA3_8 ), .B2(n216), 
        .ZN(n252) );
  AOI22_X2 U92 ( .A1(\U9/DATA8_7 ), .A2(n211), .B1(\U9/DATA7_7 ), .B2(n212), 
        .ZN(n266) );
  AOI22_X2 U93 ( .A1(\U9/DATA2_7 ), .A2(n217), .B1(\U9/DATA1_7 ), .B2(n218), 
        .ZN(n263) );
  AOI22_X2 U94 ( .A1(\U9/DATA4_7 ), .A2(n215), .B1(\U9/DATA3_7 ), .B2(n216), 
        .ZN(n264) );
  AOI22_X2 U95 ( .A1(\U9/DATA8_6 ), .A2(n211), .B1(\U9/DATA7_6 ), .B2(n212), 
        .ZN(n278) );
  AOI22_X2 U97 ( .A1(\U9/DATA2_6 ), .A2(n217), .B1(\U9/DATA1_6 ), .B2(n218), 
        .ZN(n275) );
  AOI22_X2 U98 ( .A1(\U9/DATA4_6 ), .A2(n215), .B1(\U9/DATA3_6 ), .B2(n216), 
        .ZN(n276) );
  AOI22_X2 U99 ( .A1(\U9/DATA8_5 ), .A2(n211), .B1(\U9/DATA7_5 ), .B2(n212), 
        .ZN(n290) );
  AOI22_X2 U100 ( .A1(\U9/DATA2_5 ), .A2(n217), .B1(\U9/DATA1_5 ), .B2(n218), 
        .ZN(n287) );
  AOI22_X2 U102 ( .A1(\U9/DATA4_5 ), .A2(n215), .B1(\U9/DATA3_5 ), .B2(n216), 
        .ZN(n288) );
  AOI22_X2 U104 ( .A1(\U9/DATA8_4 ), .A2(n211), .B1(\U9/DATA7_4 ), .B2(n212), 
        .ZN(n302) );
  AOI22_X2 U105 ( .A1(\U9/DATA2_4 ), .A2(n217), .B1(\U9/DATA1_4 ), .B2(n218), 
        .ZN(n299) );
  AOI22_X2 U106 ( .A1(\U9/DATA4_4 ), .A2(n215), .B1(\U9/DATA3_4 ), .B2(n216), 
        .ZN(n300) );
  AOI22_X2 U107 ( .A1(\U9/DATA8_3 ), .A2(n211), .B1(\U9/DATA7_3 ), .B2(n212), 
        .ZN(n314) );
  AOI22_X2 U109 ( .A1(\U9/DATA2_3 ), .A2(n217), .B1(\U9/DATA1_3 ), .B2(n218), 
        .ZN(n311) );
  AOI22_X2 U110 ( .A1(\U9/DATA4_3 ), .A2(n215), .B1(\U9/DATA3_3 ), .B2(n216), 
        .ZN(n312) );
  AOI22_X2 U111 ( .A1(\U9/DATA8_2 ), .A2(n211), .B1(\U9/DATA7_2 ), .B2(n212), 
        .ZN(n326) );
  AOI22_X2 U112 ( .A1(\U9/DATA2_2 ), .A2(n217), .B1(\U9/DATA1_2 ), .B2(n218), 
        .ZN(n323) );
  AOI22_X2 U114 ( .A1(\U9/DATA4_2 ), .A2(n215), .B1(\U9/DATA3_2 ), .B2(n216), 
        .ZN(n324) );
  AOI22_X2 U116 ( .A1(\U9/DATA8_1 ), .A2(n211), .B1(\U9/DATA7_1 ), .B2(n212), 
        .ZN(n338) );
  AOI22_X2 U117 ( .A1(\U9/DATA2_1 ), .A2(n217), .B1(\U9/DATA1_1 ), .B2(n218), 
        .ZN(n335) );
  AOI22_X2 U118 ( .A1(\U9/DATA4_1 ), .A2(n215), .B1(\U9/DATA3_1 ), .B2(n216), 
        .ZN(n336) );
  INV_X4 U119 ( .A(n339), .ZN(n832) );
  INV_X4 U121 ( .A(n70), .ZN(n819) );
  OAI21_X2 U122 ( .B1(n204), .B2(n205), .A(n206), .ZN(n203) );
  AOI21_X2 U123 ( .B1(n832), .B2(n837), .A(n833), .ZN(n202) );
  OAI21_X2 U124 ( .B1(n181), .B2(n182), .A(n44), .ZN(n180) );
  OAI21_X2 U126 ( .B1(n342), .B2(n343), .A(n206), .ZN(n341) );
  AOI21_X2 U129 ( .B1(n233), .B2(n234), .A(n831), .ZN(n232) );
  AOI21_X2 U130 ( .B1(n245), .B2(n246), .A(n831), .ZN(n244) );
  AOI21_X2 U131 ( .B1(n257), .B2(n258), .A(n831), .ZN(n256) );
  AOI21_X2 U132 ( .B1(n269), .B2(n270), .A(n831), .ZN(n268) );
  AOI21_X2 U136 ( .B1(n281), .B2(n282), .A(n831), .ZN(n280) );
  AOI21_X2 U137 ( .B1(n293), .B2(n294), .A(n831), .ZN(n292) );
  AOI21_X2 U138 ( .B1(n305), .B2(n306), .A(n831), .ZN(n304) );
  AOI21_X2 U140 ( .B1(n317), .B2(n318), .A(n831), .ZN(n316) );
  AOI21_X2 U146 ( .B1(n329), .B2(n330), .A(n831), .ZN(n328) );
  AOI21_X2 U149 ( .B1(n200), .B2(FoundY[0]), .A(WireY), .ZN(n70) );
  OAI21_X2 U151 ( .B1(n361), .B2(WireX), .A(DiagonalDoneX), .ZN(n339) );
  AOI22_X2 U152 ( .A1(\U8/DATA2_0 ), .A2(n55), .B1(\U8/DATA1_0 ), .B2(n56), 
        .ZN(n183) );
  AOI22_X2 U153 ( .A1(\U8/DATA10_0 ), .A2(n67), .B1(\U8/DATA9_0 ), .B2(n68), 
        .ZN(n193) );
  AOI22_X2 U154 ( .A1(\U9/DATA2_0 ), .A2(n217), .B1(\U9/DATA1_0 ), .B2(n218), 
        .ZN(n344) );
  AOI22_X2 U156 ( .A1(\U8/DATA4_0 ), .A2(n53), .B1(\U8/DATA3_0 ), .B2(n54), 
        .ZN(n184) );
  AOI22_X2 U157 ( .A1(\U8/DATA12_0 ), .A2(n65), .B1(\U8/DATA11_0 ), .B2(n66), 
        .ZN(n194) );
  AOI22_X2 U158 ( .A1(\U9/DATA4_0 ), .A2(n215), .B1(\U9/DATA3_0 ), .B2(n216), 
        .ZN(n345) );
  AOI22_X2 U159 ( .A1(\U8/DATA8_0 ), .A2(n49), .B1(\U8/DATA7_0 ), .B2(n50), 
        .ZN(n186) );
  AOI22_X2 U160 ( .A1(\U8/DATA16_0 ), .A2(n61), .B1(\U8/DATA15_0 ), .B2(n62), 
        .ZN(n196) );
  AOI22_X2 U163 ( .A1(\U9/DATA8_0 ), .A2(n211), .B1(\U9/DATA7_0 ), .B2(n212), 
        .ZN(n347) );
  AOI22_X2 U165 ( .A1(\U9/DATA16_0 ), .A2(n223), .B1(\U9/DATA15_0 ), .B2(n224), 
        .ZN(n357) );
  AOI22_X2 U166 ( .A1(\U8/DATA6_10 ), .A2(n51), .B1(\U8/DATA5_10 ), .B2(n52), 
        .ZN(n47) );
  AOI22_X2 U167 ( .A1(\U8/DATA14_10 ), .A2(n63), .B1(\U8/DATA13_10 ), .B2(n64), 
        .ZN(n59) );
  AOI22_X2 U168 ( .A1(\U8/DATA6_0 ), .A2(n51), .B1(\U8/DATA5_0 ), .B2(n52), 
        .ZN(n185) );
  AOI22_X2 U170 ( .A1(\U8/DATA14_0 ), .A2(n63), .B1(\U8/DATA13_0 ), .B2(n64), 
        .ZN(n195) );
  AOI22_X2 U171 ( .A1(\U9/DATA6_10 ), .A2(n213), .B1(\U9/DATA5_10 ), .B2(n214), 
        .ZN(n209) );
  AOI22_X2 U172 ( .A1(\U9/DATA14_10 ), .A2(n225), .B1(\U9/DATA13_10 ), .B2(
        n226), .ZN(n221) );
  AOI22_X2 U173 ( .A1(\U9/DATA6_0 ), .A2(n213), .B1(\U9/DATA5_0 ), .B2(n214), 
        .ZN(n346) );
  AOI22_X2 U175 ( .A1(\U9/DATA14_0 ), .A2(n225), .B1(\U9/DATA13_0 ), .B2(n226), 
        .ZN(n356) );
  AOI22_X2 U177 ( .A1(\U8/DATA12_9 ), .A2(n65), .B1(\U8/DATA11_9 ), .B2(n66), 
        .ZN(n77) );
  AOI22_X2 U178 ( .A1(\U8/DATA12_8 ), .A2(n65), .B1(\U8/DATA11_8 ), .B2(n66), 
        .ZN(n89) );
  AOI22_X2 U179 ( .A1(\U8/DATA12_7 ), .A2(n65), .B1(\U8/DATA11_7 ), .B2(n66), 
        .ZN(n101) );
  AOI22_X2 U180 ( .A1(\U8/DATA12_6 ), .A2(n65), .B1(\U8/DATA11_6 ), .B2(n66), 
        .ZN(n113) );
  AOI22_X2 U182 ( .A1(\U8/DATA12_5 ), .A2(n65), .B1(\U8/DATA11_5 ), .B2(n66), 
        .ZN(n125) );
  AOI22_X2 U183 ( .A1(\U8/DATA12_4 ), .A2(n65), .B1(\U8/DATA11_4 ), .B2(n66), 
        .ZN(n137) );
  AOI22_X2 U184 ( .A1(\U8/DATA12_3 ), .A2(n65), .B1(\U8/DATA11_3 ), .B2(n66), 
        .ZN(n149) );
  AOI22_X2 U185 ( .A1(\U8/DATA12_2 ), .A2(n65), .B1(\U8/DATA11_2 ), .B2(n66), 
        .ZN(n161) );
  AOI22_X2 U187 ( .A1(\U8/DATA12_1 ), .A2(n65), .B1(\U8/DATA11_1 ), .B2(n66), 
        .ZN(n173) );
  AOI22_X2 U189 ( .A1(\U8/DATA10_9 ), .A2(n67), .B1(\U8/DATA9_9 ), .B2(n68), 
        .ZN(n76) );
  AOI22_X2 U190 ( .A1(\U8/DATA10_8 ), .A2(n67), .B1(\U8/DATA9_8 ), .B2(n68), 
        .ZN(n88) );
  AOI22_X2 U191 ( .A1(\U8/DATA10_7 ), .A2(n67), .B1(\U8/DATA9_7 ), .B2(n68), 
        .ZN(n100) );
  AOI22_X2 U192 ( .A1(\U8/DATA10_6 ), .A2(n67), .B1(\U8/DATA9_6 ), .B2(n68), 
        .ZN(n112) );
  AOI22_X2 U194 ( .A1(\U8/DATA10_5 ), .A2(n67), .B1(\U8/DATA9_5 ), .B2(n68), 
        .ZN(n124) );
  AOI22_X2 U195 ( .A1(\U8/DATA10_4 ), .A2(n67), .B1(\U8/DATA9_4 ), .B2(n68), 
        .ZN(n136) );
  AOI22_X2 U196 ( .A1(\U8/DATA10_3 ), .A2(n67), .B1(\U8/DATA9_3 ), .B2(n68), 
        .ZN(n148) );
  AOI22_X2 U197 ( .A1(\U8/DATA10_2 ), .A2(n67), .B1(\U8/DATA9_2 ), .B2(n68), 
        .ZN(n160) );
  AOI22_X2 U199 ( .A1(\U8/DATA10_1 ), .A2(n67), .B1(\U8/DATA9_1 ), .B2(n68), 
        .ZN(n172) );
  AOI22_X2 U201 ( .A1(\U8/DATA16_9 ), .A2(n61), .B1(\U8/DATA15_9 ), .B2(n62), 
        .ZN(n79) );
  AOI22_X2 U202 ( .A1(\U8/DATA16_8 ), .A2(n61), .B1(\U8/DATA15_8 ), .B2(n62), 
        .ZN(n91) );
  AOI22_X2 U203 ( .A1(\U8/DATA16_7 ), .A2(n61), .B1(\U8/DATA15_7 ), .B2(n62), 
        .ZN(n103) );
  AOI22_X2 U204 ( .A1(\U8/DATA16_6 ), .A2(n61), .B1(\U8/DATA15_6 ), .B2(n62), 
        .ZN(n115) );
  AOI22_X2 U206 ( .A1(\U8/DATA16_5 ), .A2(n61), .B1(\U8/DATA15_5 ), .B2(n62), 
        .ZN(n127) );
  AOI22_X2 U207 ( .A1(\U8/DATA16_4 ), .A2(n61), .B1(\U8/DATA15_4 ), .B2(n62), 
        .ZN(n139) );
  AOI22_X2 U208 ( .A1(\U8/DATA16_3 ), .A2(n61), .B1(\U8/DATA15_3 ), .B2(n62), 
        .ZN(n151) );
  AOI22_X2 U209 ( .A1(\U8/DATA16_2 ), .A2(n61), .B1(\U8/DATA15_2 ), .B2(n62), 
        .ZN(n163) );
  AOI22_X2 U211 ( .A1(\U8/DATA16_1 ), .A2(n61), .B1(\U8/DATA15_1 ), .B2(n62), 
        .ZN(n175) );
  AOI22_X2 U213 ( .A1(\U9/DATA16_9 ), .A2(n223), .B1(\U9/DATA15_9 ), .B2(n224), 
        .ZN(n238) );
  AOI22_X2 U214 ( .A1(\U9/DATA16_8 ), .A2(n223), .B1(\U9/DATA15_8 ), .B2(n224), 
        .ZN(n250) );
  AOI22_X2 U215 ( .A1(\U9/DATA16_7 ), .A2(n223), .B1(\U9/DATA15_7 ), .B2(n224), 
        .ZN(n262) );
  AOI22_X2 U216 ( .A1(\U9/DATA16_6 ), .A2(n223), .B1(\U9/DATA15_6 ), .B2(n224), 
        .ZN(n274) );
  AOI22_X2 U218 ( .A1(\U9/DATA16_5 ), .A2(n223), .B1(\U9/DATA15_5 ), .B2(n224), 
        .ZN(n286) );
  AOI22_X2 U219 ( .A1(\U9/DATA16_4 ), .A2(n223), .B1(\U9/DATA15_4 ), .B2(n224), 
        .ZN(n298) );
  AOI22_X2 U220 ( .A1(\U9/DATA16_3 ), .A2(n223), .B1(\U9/DATA15_3 ), .B2(n224), 
        .ZN(n310) );
  AOI22_X2 U221 ( .A1(\U9/DATA16_2 ), .A2(n223), .B1(\U9/DATA15_2 ), .B2(n224), 
        .ZN(n322) );
  AOI22_X2 U223 ( .A1(\U9/DATA16_1 ), .A2(n223), .B1(\U9/DATA15_1 ), .B2(n224), 
        .ZN(n334) );
  AOI22_X2 U225 ( .A1(\U8/DATA6_9 ), .A2(n51), .B1(\U8/DATA5_9 ), .B2(n52), 
        .ZN(n82) );
  AOI22_X2 U226 ( .A1(\U8/DATA14_9 ), .A2(n63), .B1(\U8/DATA13_9 ), .B2(n64), 
        .ZN(n78) );
  AOI22_X2 U227 ( .A1(\U8/DATA6_8 ), .A2(n51), .B1(\U8/DATA5_8 ), .B2(n52), 
        .ZN(n94) );
  AOI22_X2 U228 ( .A1(\U8/DATA14_8 ), .A2(n63), .B1(\U8/DATA13_8 ), .B2(n64), 
        .ZN(n90) );
  AOI22_X2 U230 ( .A1(\U8/DATA6_7 ), .A2(n51), .B1(\U8/DATA5_7 ), .B2(n52), 
        .ZN(n106) );
  AOI22_X2 U231 ( .A1(\U8/DATA14_7 ), .A2(n63), .B1(\U8/DATA13_7 ), .B2(n64), 
        .ZN(n102) );
  AOI22_X2 U232 ( .A1(\U8/DATA6_6 ), .A2(n51), .B1(\U8/DATA5_6 ), .B2(n52), 
        .ZN(n118) );
  AOI22_X2 U233 ( .A1(\U8/DATA14_6 ), .A2(n63), .B1(\U8/DATA13_6 ), .B2(n64), 
        .ZN(n114) );
  AOI22_X2 U235 ( .A1(\U8/DATA6_5 ), .A2(n51), .B1(\U8/DATA5_5 ), .B2(n52), 
        .ZN(n130) );
  AOI22_X2 U237 ( .A1(\U8/DATA14_5 ), .A2(n63), .B1(\U8/DATA13_5 ), .B2(n64), 
        .ZN(n126) );
  AOI22_X2 U238 ( .A1(\U8/DATA6_4 ), .A2(n51), .B1(\U8/DATA5_4 ), .B2(n52), 
        .ZN(n142) );
  AOI22_X2 U239 ( .A1(\U8/DATA14_4 ), .A2(n63), .B1(\U8/DATA13_4 ), .B2(n64), 
        .ZN(n138) );
  AOI22_X2 U240 ( .A1(\U8/DATA6_3 ), .A2(n51), .B1(\U8/DATA5_3 ), .B2(n52), 
        .ZN(n154) );
  AOI22_X2 U242 ( .A1(\U8/DATA14_3 ), .A2(n63), .B1(\U8/DATA13_3 ), .B2(n64), 
        .ZN(n150) );
  AOI22_X2 U243 ( .A1(\U8/DATA6_2 ), .A2(n51), .B1(\U8/DATA5_2 ), .B2(n52), 
        .ZN(n166) );
  AOI22_X2 U244 ( .A1(\U8/DATA14_2 ), .A2(n63), .B1(\U8/DATA13_2 ), .B2(n64), 
        .ZN(n162) );
  AOI22_X2 U245 ( .A1(\U8/DATA6_1 ), .A2(n51), .B1(\U8/DATA5_1 ), .B2(n52), 
        .ZN(n178) );
  AOI22_X2 U247 ( .A1(\U8/DATA14_1 ), .A2(n63), .B1(\U8/DATA13_1 ), .B2(n64), 
        .ZN(n174) );
  AOI22_X2 U249 ( .A1(\U9/DATA6_9 ), .A2(n213), .B1(\U9/DATA5_9 ), .B2(n214), 
        .ZN(n241) );
  AOI22_X2 U250 ( .A1(\U9/DATA14_9 ), .A2(n225), .B1(\U9/DATA13_9 ), .B2(n226), 
        .ZN(n237) );
  AOI22_X2 U251 ( .A1(\U9/DATA6_8 ), .A2(n213), .B1(\U9/DATA5_8 ), .B2(n214), 
        .ZN(n253) );
  AOI22_X2 U252 ( .A1(\U9/DATA14_8 ), .A2(n225), .B1(\U9/DATA13_8 ), .B2(n226), 
        .ZN(n249) );
  AOI22_X2 U254 ( .A1(\U9/DATA6_7 ), .A2(n213), .B1(\U9/DATA5_7 ), .B2(n214), 
        .ZN(n265) );
  AOI22_X2 U255 ( .A1(\U9/DATA14_7 ), .A2(n225), .B1(\U9/DATA13_7 ), .B2(n226), 
        .ZN(n261) );
  AOI22_X2 U256 ( .A1(\U9/DATA6_6 ), .A2(n213), .B1(\U9/DATA5_6 ), .B2(n214), 
        .ZN(n277) );
  AOI22_X2 U257 ( .A1(\U9/DATA14_6 ), .A2(n225), .B1(\U9/DATA13_6 ), .B2(n226), 
        .ZN(n273) );
  AOI22_X2 U259 ( .A1(\U9/DATA6_5 ), .A2(n213), .B1(\U9/DATA5_5 ), .B2(n214), 
        .ZN(n289) );
  AOI22_X2 U261 ( .A1(\U9/DATA14_5 ), .A2(n225), .B1(\U9/DATA13_5 ), .B2(n226), 
        .ZN(n285) );
  AOI22_X2 U262 ( .A1(\U9/DATA6_4 ), .A2(n213), .B1(\U9/DATA5_4 ), .B2(n214), 
        .ZN(n301) );
  AOI22_X2 U263 ( .A1(\U9/DATA14_4 ), .A2(n225), .B1(\U9/DATA13_4 ), .B2(n226), 
        .ZN(n297) );
  AOI22_X2 U264 ( .A1(\U9/DATA6_3 ), .A2(n213), .B1(\U9/DATA5_3 ), .B2(n214), 
        .ZN(n313) );
  AOI22_X2 U266 ( .A1(\U9/DATA14_3 ), .A2(n225), .B1(\U9/DATA13_3 ), .B2(n226), 
        .ZN(n309) );
  AOI22_X2 U267 ( .A1(\U9/DATA6_2 ), .A2(n213), .B1(\U9/DATA5_2 ), .B2(n214), 
        .ZN(n325) );
  AOI22_X2 U268 ( .A1(\U9/DATA14_2 ), .A2(n225), .B1(\U9/DATA13_2 ), .B2(n226), 
        .ZN(n321) );
  AOI22_X2 U269 ( .A1(\U9/DATA6_1 ), .A2(n213), .B1(\U9/DATA5_1 ), .B2(n214), 
        .ZN(n337) );
  AOI22_X2 U271 ( .A1(\U9/DATA14_1 ), .A2(n225), .B1(\U9/DATA13_1 ), .B2(n226), 
        .ZN(n333) );
  OAI211_X2 U274 ( .C1(n821), .C2(n13), .A(n40), .B(n41), .ZN(n362) );
  OAI21_X2 U275 ( .B1(n42), .B2(n43), .A(n44), .ZN(n41) );
  AOI21_X2 U276 ( .B1(n74), .B2(n75), .A(n818), .ZN(n73) );
  AOI21_X2 U277 ( .B1(n86), .B2(n87), .A(n818), .ZN(n85) );
  AOI21_X2 U281 ( .B1(n98), .B2(n99), .A(n818), .ZN(n97) );
  AOI21_X2 U282 ( .B1(n110), .B2(n111), .A(n818), .ZN(n109) );
  AOI21_X2 U283 ( .B1(n122), .B2(n123), .A(n818), .ZN(n121) );
  AOI21_X2 U285 ( .B1(n134), .B2(n135), .A(n818), .ZN(n133) );
  AOI21_X2 U291 ( .B1(n146), .B2(n147), .A(n818), .ZN(n145) );
  AOI21_X2 U293 ( .B1(n158), .B2(n159), .A(n818), .ZN(n157) );
  AOI21_X2 U294 ( .B1(n170), .B2(n171), .A(n818), .ZN(n169) );
  AND2_X4 U295 ( .A1(n353), .A2(n359), .ZN(n229) );
  AND2_X4 U296 ( .A1(n353), .A2(n358), .ZN(n230) );
  AND2_X4 U297 ( .A1(n352), .A2(n359), .ZN(n227) );
  AND2_X4 U298 ( .A1(n352), .A2(n358), .ZN(n228) );
  AND2_X4 U299 ( .A1(n351), .A2(n359), .ZN(n225) );
  AND2_X4 U300 ( .A1(n351), .A2(n358), .ZN(n226) );
  AND2_X4 U301 ( .A1(n349), .A2(n359), .ZN(n223) );
  AND2_X4 U302 ( .A1(n358), .A2(n349), .ZN(n224) );
  AND2_X4 U303 ( .A1(n350), .A2(n353), .ZN(n217) );
  AND2_X4 U304 ( .A1(n348), .A2(n353), .ZN(n218) );
  AND2_X4 U305 ( .A1(n350), .A2(n352), .ZN(n215) );
  AND2_X4 U306 ( .A1(n348), .A2(n352), .ZN(n216) );
  AND2_X4 U307 ( .A1(n350), .A2(n351), .ZN(n213) );
  AND2_X4 U308 ( .A1(n348), .A2(n351), .ZN(n214) );
  AND2_X4 U309 ( .A1(n350), .A2(n349), .ZN(n211) );
  AND2_X4 U310 ( .A1(n348), .A2(n349), .ZN(n212) );
  AND2_X4 U311 ( .A1(n192), .A2(n198), .ZN(n67) );
  AND2_X4 U312 ( .A1(n192), .A2(n197), .ZN(n68) );
  AND2_X4 U313 ( .A1(n191), .A2(n198), .ZN(n65) );
  AND2_X4 U314 ( .A1(n191), .A2(n197), .ZN(n66) );
  AND2_X4 U315 ( .A1(n190), .A2(n198), .ZN(n63) );
  AND2_X4 U316 ( .A1(n190), .A2(n197), .ZN(n64) );
  AND2_X4 U317 ( .A1(n188), .A2(n198), .ZN(n61) );
  AND2_X4 U318 ( .A1(n197), .A2(n188), .ZN(n62) );
  AND2_X4 U319 ( .A1(n189), .A2(n192), .ZN(n55) );
  AND2_X4 U320 ( .A1(n187), .A2(n192), .ZN(n56) );
  AND2_X4 U321 ( .A1(n189), .A2(n191), .ZN(n53) );
  AND2_X4 U322 ( .A1(n187), .A2(n191), .ZN(n54) );
  AND2_X4 U323 ( .A1(n189), .A2(n190), .ZN(n51) );
  AND2_X4 U324 ( .A1(n187), .A2(n190), .ZN(n52) );
  AND2_X4 U325 ( .A1(n189), .A2(n188), .ZN(n49) );
  AND2_X4 U326 ( .A1(n187), .A2(n188), .ZN(n50) );
  INV_X4 U327 ( .A(n72), .ZN(n809) );
  INV_X4 U328 ( .A(n84), .ZN(n810) );
  INV_X4 U329 ( .A(n96), .ZN(n811) );
  INV_X4 U330 ( .A(n108), .ZN(n812) );
  INV_X4 U331 ( .A(n120), .ZN(n813) );
  INV_X4 U332 ( .A(n132), .ZN(n814) );
  INV_X4 U333 ( .A(n144), .ZN(n815) );
  INV_X4 U334 ( .A(n156), .ZN(n816) );
  INV_X4 U335 ( .A(n168), .ZN(n817) );
  INV_X4 U336 ( .A(n44), .ZN(n818) );
  INV_X4 U337 ( .A(n71), .ZN(n820) );
  INV_X4 U339 ( .A(n69), .ZN(n821) );
  INV_X4 U340 ( .A(n231), .ZN(n822) );
  INV_X4 U342 ( .A(n243), .ZN(n823) );
  INV_X4 U343 ( .A(n255), .ZN(n824) );
  INV_X4 U344 ( .A(n267), .ZN(n825) );
  INV_X4 U345 ( .A(n279), .ZN(n826) );
  INV_X4 U346 ( .A(n291), .ZN(n827) );
  INV_X4 U347 ( .A(n303), .ZN(n828) );
  INV_X4 U348 ( .A(n315), .ZN(n829) );
  INV_X4 U349 ( .A(n327), .ZN(n830) );
  INV_X4 U350 ( .A(n206), .ZN(n831) );
  INV_X4 U351 ( .A(n340), .ZN(n833) );
  INV_X4 U352 ( .A(FoundX[0]), .ZN(n834) );
  INV_X4 U353 ( .A(DiagonalDoneX), .ZN(n835) );
  INV_X4 U354 ( .A(DiagonalDoneY), .ZN(n836) );
  INV_X4 U355 ( .A(\add_87/carry[10] ), .ZN(n837) );
  INV_X4 U357 ( .A(X[3]), .ZN(n838) );
  INV_X4 U358 ( .A(X[1]), .ZN(n839) );
  INV_X4 U360 ( .A(X[0]), .ZN(n840) );
  INV_X4 U361 ( .A(Y[3]), .ZN(n841) );
  INV_X4 U362 ( .A(Y[1]), .ZN(n842) );
  INV_X4 U363 ( .A(Y[0]), .ZN(n843) );
endmodule


module MainArbiter_1 ( reset, clock, EnableChange, Update_1Req1, Update_1Req2, 
        Update_2Req1, Update_2Req2, Row1, Row2, OutputReq1, OutputReq2, 
        Output_1Row1, Output_1Row2, Output_2Row1, Output_2Row2, FlagX, FlagY, 
        DiagonalDoneX, DiagonalDoneY, WE, PosDX, PaddedRow, WriteReq, WriteBus, 
        NewDiagonalX, NewDiagonalY, NewElement, ArbiterElement, ArbiterPos, 
        OutputPaddedRow, PosDY, PosRowX, PosRowY, ComputeReq, OutputCompute, 
        CompStart, EOC_Flag );
  input [10:0] Update_1Req1;
  input [10:0] Update_1Req2;
  input [10:0] Update_2Req1;
  input [10:0] Update_2Req2;
  input [255:0] Row1;
  input [255:0] Row2;
  output [10:0] OutputReq1;
  output [10:0] OutputReq2;
  output [255:0] Output_1Row1;
  output [255:0] Output_1Row2;
  output [255:0] Output_2Row1;
  output [255:0] Output_2Row2;
  input [12:0] PosDX;
  input [255:0] PaddedRow;
  output [10:0] WriteReq;
  output [255:0] WriteBus;
  input [47:0] NewDiagonalX;
  input [47:0] NewDiagonalY;
  input [47:0] NewElement;
  output [47:0] ArbiterElement;
  output [12:0] ArbiterPos;
  output [255:0] OutputPaddedRow;
  input [12:0] PosDY;
  input [12:0] PosRowX;
  input [12:0] PosRowY;
  input [10:0] ComputeReq;
  output [255:0] OutputCompute;
  input reset, clock, EnableChange, DiagonalDoneX, DiagonalDoneY, EOC_Flag;
  output FlagX, FlagY, WE, CompStart;
  wire   n1830, n1828, \U3/U1/Z_0 , \U3/U2/Z_0 , \U3/U3/Z_0 , \U3/U3/Z_1 ,
         \U3/U3/Z_2 , \U3/U3/Z_3 , \U3/U3/Z_4 , \U3/U3/Z_5 , \U3/U3/Z_6 ,
         \U3/U3/Z_7 , \U3/U3/Z_8 , \U3/U3/Z_9 , \U3/U3/Z_10 , \U3/U3/DATA2_0 ,
         \U3/U3/DATA2_1 , \U3/U3/DATA2_2 , \U3/U3/DATA2_3 , \U3/U3/DATA2_4 ,
         \U3/U3/DATA2_5 , \U3/U3/DATA2_6 , \U3/U3/DATA2_7 , \U3/U3/DATA2_8 ,
         \U3/U3/DATA2_9 , \U3/U3/DATA2_10 , \U3/U3/DATA1_0 , \U3/U3/DATA1_1 ,
         \U3/U3/DATA1_2 , \U3/U3/DATA1_3 , \U3/U3/DATA1_4 , \U3/U3/DATA1_5 ,
         \U3/U3/DATA1_6 , \U3/U3/DATA1_7 , \U3/U3/DATA1_8 , \U3/U3/DATA1_9 ,
         \U3/U3/DATA1_10 , \U3/U4/DATA2_0 , \U3/U5/Z_0 , \U3/U5/Z_1 ,
         \U3/U5/Z_2 , \U3/U5/Z_3 , \U3/U5/Z_4 , \U3/U5/Z_5 , \U3/U5/Z_6 ,
         \U3/U5/Z_7 , \U3/U5/Z_8 , \U3/U5/Z_9 , \U3/U5/Z_10 , \U3/U5/Z_11 ,
         \U3/U5/Z_12 , \U3/U5/Z_13 , \U3/U5/Z_14 , \U3/U5/Z_15 , \U3/U5/Z_16 ,
         \U3/U5/Z_17 , \U3/U5/Z_18 , \U3/U5/Z_19 , \U3/U5/Z_20 , \U3/U5/Z_21 ,
         \U3/U5/Z_22 , \U3/U5/Z_23 , \U3/U5/Z_24 , \U3/U5/Z_25 , \U3/U5/Z_26 ,
         \U3/U5/Z_27 , \U3/U5/Z_28 , \U3/U5/Z_29 , \U3/U5/Z_30 , \U3/U5/Z_31 ,
         \U3/U5/Z_32 , \U3/U5/Z_33 , \U3/U5/Z_34 , \U3/U5/Z_35 , \U3/U5/Z_36 ,
         \U3/U5/Z_37 , \U3/U5/Z_38 , \U3/U5/Z_39 , \U3/U5/Z_40 , \U3/U5/Z_41 ,
         \U3/U5/Z_42 , \U3/U5/Z_43 , \U3/U5/Z_44 , \U3/U5/Z_45 , \U3/U5/Z_46 ,
         \U3/U5/Z_47 , \U3/U5/DATA3_0 , \U3/U5/DATA3_1 , \U3/U5/DATA3_2 ,
         \U3/U5/DATA3_3 , \U3/U5/DATA3_4 , \U3/U5/DATA3_5 , \U3/U5/DATA3_6 ,
         \U3/U5/DATA3_7 , \U3/U5/DATA3_8 , \U3/U5/DATA3_9 , \U3/U5/DATA3_10 ,
         \U3/U5/DATA3_11 , \U3/U5/DATA3_12 , \U3/U5/DATA3_13 ,
         \U3/U5/DATA3_14 , \U3/U5/DATA3_15 , \U3/U5/DATA3_16 ,
         \U3/U5/DATA3_17 , \U3/U5/DATA3_18 , \U3/U5/DATA3_19 ,
         \U3/U5/DATA3_20 , \U3/U5/DATA3_21 , \U3/U5/DATA3_22 ,
         \U3/U5/DATA3_23 , \U3/U5/DATA3_24 , \U3/U5/DATA3_25 ,
         \U3/U5/DATA3_26 , \U3/U5/DATA3_27 , \U3/U5/DATA3_28 ,
         \U3/U5/DATA3_29 , \U3/U5/DATA3_30 , \U3/U5/DATA3_31 ,
         \U3/U5/DATA3_32 , \U3/U5/DATA3_33 , \U3/U5/DATA3_34 ,
         \U3/U5/DATA3_35 , \U3/U5/DATA3_36 , \U3/U5/DATA3_37 ,
         \U3/U5/DATA3_38 , \U3/U5/DATA3_39 , \U3/U5/DATA3_40 ,
         \U3/U5/DATA3_41 , \U3/U5/DATA3_42 , \U3/U5/DATA3_43 ,
         \U3/U5/DATA3_44 , \U3/U5/DATA3_45 , \U3/U5/DATA3_46 ,
         \U3/U5/DATA3_47 , \U3/U5/DATA2_0 , \U3/U5/DATA2_1 , \U3/U5/DATA2_2 ,
         \U3/U5/DATA2_3 , \U3/U5/DATA2_4 , \U3/U5/DATA2_5 , \U3/U5/DATA2_6 ,
         \U3/U5/DATA2_7 , \U3/U5/DATA2_8 , \U3/U5/DATA2_9 , \U3/U5/DATA2_10 ,
         \U3/U5/DATA2_11 , \U3/U5/DATA2_12 , \U3/U5/DATA2_13 ,
         \U3/U5/DATA2_14 , \U3/U5/DATA2_15 , \U3/U5/DATA2_16 ,
         \U3/U5/DATA2_17 , \U3/U5/DATA2_18 , \U3/U5/DATA2_19 ,
         \U3/U5/DATA2_20 , \U3/U5/DATA2_21 , \U3/U5/DATA2_22 ,
         \U3/U5/DATA2_23 , \U3/U5/DATA2_24 , \U3/U5/DATA2_25 ,
         \U3/U5/DATA2_26 , \U3/U5/DATA2_27 , \U3/U5/DATA2_28 ,
         \U3/U5/DATA2_29 , \U3/U5/DATA2_30 , \U3/U5/DATA2_31 ,
         \U3/U5/DATA2_32 , \U3/U5/DATA2_33 , \U3/U5/DATA2_34 ,
         \U3/U5/DATA2_35 , \U3/U5/DATA2_36 , \U3/U5/DATA2_37 ,
         \U3/U5/DATA2_38 , \U3/U5/DATA2_39 , \U3/U5/DATA2_40 ,
         \U3/U5/DATA2_41 , \U3/U5/DATA2_42 , \U3/U5/DATA2_43 ,
         \U3/U5/DATA2_44 , \U3/U5/DATA2_45 , \U3/U5/DATA2_46 ,
         \U3/U5/DATA2_47 , \U3/U5/DATA1_0 , \U3/U5/DATA1_1 , \U3/U5/DATA1_2 ,
         \U3/U5/DATA1_3 , \U3/U5/DATA1_4 , \U3/U5/DATA1_5 , \U3/U5/DATA1_6 ,
         \U3/U5/DATA1_7 , \U3/U5/DATA1_8 , \U3/U5/DATA1_9 , \U3/U5/DATA1_10 ,
         \U3/U5/DATA1_11 , \U3/U5/DATA1_12 , \U3/U5/DATA1_13 ,
         \U3/U5/DATA1_14 , \U3/U5/DATA1_15 , \U3/U5/DATA1_16 ,
         \U3/U5/DATA1_17 , \U3/U5/DATA1_18 , \U3/U5/DATA1_19 ,
         \U3/U5/DATA1_20 , \U3/U5/DATA1_21 , \U3/U5/DATA1_22 ,
         \U3/U5/DATA1_23 , \U3/U5/DATA1_24 , \U3/U5/DATA1_25 ,
         \U3/U5/DATA1_26 , \U3/U5/DATA1_27 , \U3/U5/DATA1_28 ,
         \U3/U5/DATA1_29 , \U3/U5/DATA1_30 , \U3/U5/DATA1_31 ,
         \U3/U5/DATA1_32 , \U3/U5/DATA1_33 , \U3/U5/DATA1_34 ,
         \U3/U5/DATA1_35 , \U3/U5/DATA1_36 , \U3/U5/DATA1_37 ,
         \U3/U5/DATA1_38 , \U3/U5/DATA1_39 , \U3/U5/DATA1_40 ,
         \U3/U5/DATA1_41 , \U3/U5/DATA1_42 , \U3/U5/DATA1_43 ,
         \U3/U5/DATA1_44 , \U3/U5/DATA1_45 , \U3/U5/DATA1_46 ,
         \U3/U5/DATA1_47 , \U3/U7/Z_0 , \U3/U7/Z_1 , \U3/U7/Z_2 , \U3/U7/Z_3 ,
         \U3/U7/Z_4 , \U3/U7/Z_5 , \U3/U7/Z_6 , \U3/U7/Z_7 , \U3/U7/Z_8 ,
         \U3/U7/Z_9 , \U3/U7/Z_10 , \U3/U7/DATA7_0 , \U3/U7/DATA7_1 ,
         \U3/U7/DATA7_2 , \U3/U7/DATA7_3 , \U3/U7/DATA7_4 , \U3/U7/DATA7_5 ,
         \U3/U7/DATA7_6 , \U3/U7/DATA7_7 , \U3/U7/DATA7_8 , \U3/U7/DATA7_9 ,
         \U3/U7/DATA7_10 , \U3/U7/DATA6_0 , \U3/U7/DATA6_1 , \U3/U7/DATA6_2 ,
         \U3/U7/DATA6_3 , \U3/U7/DATA6_4 , \U3/U7/DATA6_5 , \U3/U7/DATA6_6 ,
         \U3/U7/DATA6_7 , \U3/U7/DATA6_8 , \U3/U7/DATA6_9 , \U3/U7/DATA6_10 ,
         \U3/U7/DATA5_0 , \U3/U7/DATA5_1 , \U3/U7/DATA5_2 , \U3/U7/DATA5_3 ,
         \U3/U7/DATA5_4 , \U3/U7/DATA5_5 , \U3/U7/DATA5_6 , \U3/U7/DATA5_7 ,
         \U3/U7/DATA5_8 , \U3/U7/DATA5_9 , \U3/U7/DATA5_10 , \U3/U7/DATA4_0 ,
         \U3/U7/DATA4_1 , \U3/U7/DATA4_2 , \U3/U7/DATA4_3 , \U3/U7/DATA4_4 ,
         \U3/U7/DATA4_5 , \U3/U7/DATA4_6 , \U3/U7/DATA4_7 , \U3/U7/DATA4_8 ,
         \U3/U7/DATA4_9 , \U3/U7/DATA4_10 , \U3/U7/DATA3_0 , \U3/U7/DATA3_1 ,
         \U3/U7/DATA3_2 , \U3/U7/DATA3_3 , \U3/U7/DATA3_4 , \U3/U7/DATA3_5 ,
         \U3/U7/DATA3_6 , \U3/U7/DATA3_7 , \U3/U7/DATA3_8 , \U3/U7/DATA3_9 ,
         \U3/U7/DATA3_10 , \U3/U7/DATA2_0 , \U3/U7/DATA2_1 , \U3/U7/DATA2_2 ,
         \U3/U7/DATA2_3 , \U3/U7/DATA2_4 , \U3/U7/DATA2_5 , \U3/U7/DATA2_6 ,
         \U3/U7/DATA2_7 , \U3/U7/DATA2_8 , \U3/U7/DATA2_9 , \U3/U7/DATA2_10 ,
         \U3/U7/DATA1_0 , \U3/U7/DATA1_1 , \U3/U7/DATA1_2 , \U3/U7/DATA1_3 ,
         \U3/U7/DATA1_4 , \U3/U7/DATA1_5 , \U3/U7/DATA1_6 , \U3/U7/DATA1_7 ,
         \U3/U7/DATA1_8 , \U3/U7/DATA1_9 , \U3/U7/DATA1_10 , \U3/U8/Z_0 ,
         \U3/U8/Z_1 , \U3/U8/DATA4_0 , \U3/U8/DATA4_1 , \U3/U8/DATA3_0 ,
         \U3/U8/DATA3_1 , \U3/U8/DATA2_0 , \U3/U8/DATA2_1 , \U3/U8/DATA1_0 ,
         \U3/U8/DATA1_1 , \U3/U9/Z_0 , \U3/U9/Z_1 , \U3/U9/Z_2 , \U3/U9/Z_3 ,
         \U3/U9/Z_4 , \U3/U9/Z_5 , \U3/U9/Z_6 , \U3/U9/Z_7 , \U3/U9/Z_8 ,
         \U3/U9/Z_9 , \U3/U9/Z_10 , \U3/U10/DATA3_0 , \U3/U10/DATA1_0 ,
         \U4/Z_0 , \U4/Z_1 , \U4/Z_3 , n8, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n2958, n2959,
         n2960, n2961, n2962, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802;
  assign WE = \U3/U1/Z_0 ;
  assign FlagY = \U3/U2/Z_0 ;
  assign OutputReq2[0] = \U3/U3/Z_0 ;
  assign OutputReq2[1] = \U3/U3/Z_1 ;
  assign OutputReq2[2] = \U3/U3/Z_2 ;
  assign OutputReq2[3] = \U3/U3/Z_3 ;
  assign OutputReq2[4] = \U3/U3/Z_4 ;
  assign OutputReq2[5] = \U3/U3/Z_5 ;
  assign OutputReq2[6] = \U3/U3/Z_6 ;
  assign OutputReq2[7] = \U3/U3/Z_7 ;
  assign OutputReq2[8] = \U3/U3/Z_8 ;
  assign OutputReq2[9] = \U3/U3/Z_9 ;
  assign OutputReq2[10] = \U3/U3/Z_10 ;
  assign \U3/U3/DATA2_0  = Update_2Req2[0];
  assign \U3/U3/DATA2_1  = Update_2Req2[1];
  assign \U3/U3/DATA2_2  = Update_2Req2[2];
  assign \U3/U3/DATA2_3  = Update_2Req2[3];
  assign \U3/U3/DATA2_4  = Update_2Req2[4];
  assign \U3/U3/DATA2_5  = Update_2Req2[5];
  assign \U3/U3/DATA2_6  = Update_2Req2[6];
  assign \U3/U3/DATA2_7  = Update_2Req2[7];
  assign \U3/U3/DATA2_8  = Update_2Req2[8];
  assign \U3/U3/DATA2_9  = Update_2Req2[9];
  assign \U3/U3/DATA2_10  = Update_2Req2[10];
  assign \U3/U3/DATA1_0  = Update_1Req2[0];
  assign \U3/U3/DATA1_1  = Update_1Req2[1];
  assign \U3/U3/DATA1_2  = Update_1Req2[2];
  assign \U3/U3/DATA1_3  = Update_1Req2[3];
  assign \U3/U3/DATA1_4  = Update_1Req2[4];
  assign \U3/U3/DATA1_5  = Update_1Req2[5];
  assign \U3/U3/DATA1_6  = Update_1Req2[6];
  assign \U3/U3/DATA1_7  = Update_1Req2[7];
  assign \U3/U3/DATA1_8  = Update_1Req2[8];
  assign \U3/U3/DATA1_9  = Update_1Req2[9];
  assign \U3/U3/DATA1_10  = Update_1Req2[10];
  assign \U3/U4/DATA2_0  = DiagonalDoneY;
  assign ArbiterElement[0] = \U3/U5/Z_0 ;
  assign ArbiterElement[1] = \U3/U5/Z_1 ;
  assign ArbiterElement[2] = \U3/U5/Z_2 ;
  assign ArbiterElement[3] = \U3/U5/Z_3 ;
  assign ArbiterElement[4] = \U3/U5/Z_4 ;
  assign ArbiterElement[5] = \U3/U5/Z_5 ;
  assign ArbiterElement[6] = \U3/U5/Z_6 ;
  assign ArbiterElement[7] = \U3/U5/Z_7 ;
  assign ArbiterElement[8] = \U3/U5/Z_8 ;
  assign ArbiterElement[9] = \U3/U5/Z_9 ;
  assign ArbiterElement[10] = \U3/U5/Z_10 ;
  assign ArbiterElement[11] = \U3/U5/Z_11 ;
  assign ArbiterElement[12] = \U3/U5/Z_12 ;
  assign ArbiterElement[13] = \U3/U5/Z_13 ;
  assign ArbiterElement[14] = \U3/U5/Z_14 ;
  assign ArbiterElement[15] = \U3/U5/Z_15 ;
  assign ArbiterElement[16] = \U3/U5/Z_16 ;
  assign ArbiterElement[17] = \U3/U5/Z_17 ;
  assign ArbiterElement[18] = \U3/U5/Z_18 ;
  assign ArbiterElement[19] = \U3/U5/Z_19 ;
  assign ArbiterElement[20] = \U3/U5/Z_20 ;
  assign ArbiterElement[21] = \U3/U5/Z_21 ;
  assign ArbiterElement[22] = \U3/U5/Z_22 ;
  assign ArbiterElement[23] = \U3/U5/Z_23 ;
  assign ArbiterElement[24] = \U3/U5/Z_24 ;
  assign ArbiterElement[25] = \U3/U5/Z_25 ;
  assign ArbiterElement[26] = \U3/U5/Z_26 ;
  assign ArbiterElement[27] = \U3/U5/Z_27 ;
  assign ArbiterElement[28] = \U3/U5/Z_28 ;
  assign ArbiterElement[29] = \U3/U5/Z_29 ;
  assign ArbiterElement[30] = \U3/U5/Z_30 ;
  assign ArbiterElement[31] = \U3/U5/Z_31 ;
  assign ArbiterElement[32] = \U3/U5/Z_32 ;
  assign ArbiterElement[33] = \U3/U5/Z_33 ;
  assign ArbiterElement[34] = \U3/U5/Z_34 ;
  assign ArbiterElement[35] = \U3/U5/Z_35 ;
  assign ArbiterElement[36] = \U3/U5/Z_36 ;
  assign ArbiterElement[37] = \U3/U5/Z_37 ;
  assign ArbiterElement[38] = \U3/U5/Z_38 ;
  assign ArbiterElement[39] = \U3/U5/Z_39 ;
  assign ArbiterElement[40] = \U3/U5/Z_40 ;
  assign ArbiterElement[41] = \U3/U5/Z_41 ;
  assign ArbiterElement[42] = \U3/U5/Z_42 ;
  assign ArbiterElement[43] = \U3/U5/Z_43 ;
  assign ArbiterElement[44] = \U3/U5/Z_44 ;
  assign ArbiterElement[45] = \U3/U5/Z_45 ;
  assign ArbiterElement[46] = \U3/U5/Z_46 ;
  assign ArbiterElement[47] = \U3/U5/Z_47 ;
  assign \U3/U5/DATA3_0  = NewElement[0];
  assign \U3/U5/DATA3_1  = NewElement[1];
  assign \U3/U5/DATA3_2  = NewElement[2];
  assign \U3/U5/DATA3_3  = NewElement[3];
  assign \U3/U5/DATA3_4  = NewElement[4];
  assign \U3/U5/DATA3_5  = NewElement[5];
  assign \U3/U5/DATA3_6  = NewElement[6];
  assign \U3/U5/DATA3_7  = NewElement[7];
  assign \U3/U5/DATA3_8  = NewElement[8];
  assign \U3/U5/DATA3_9  = NewElement[9];
  assign \U3/U5/DATA3_10  = NewElement[10];
  assign \U3/U5/DATA3_11  = NewElement[11];
  assign \U3/U5/DATA3_12  = NewElement[12];
  assign \U3/U5/DATA3_13  = NewElement[13];
  assign \U3/U5/DATA3_14  = NewElement[14];
  assign \U3/U5/DATA3_15  = NewElement[15];
  assign \U3/U5/DATA3_16  = NewElement[16];
  assign \U3/U5/DATA3_17  = NewElement[17];
  assign \U3/U5/DATA3_18  = NewElement[18];
  assign \U3/U5/DATA3_19  = NewElement[19];
  assign \U3/U5/DATA3_20  = NewElement[20];
  assign \U3/U5/DATA3_21  = NewElement[21];
  assign \U3/U5/DATA3_22  = NewElement[22];
  assign \U3/U5/DATA3_23  = NewElement[23];
  assign \U3/U5/DATA3_24  = NewElement[24];
  assign \U3/U5/DATA3_25  = NewElement[25];
  assign \U3/U5/DATA3_26  = NewElement[26];
  assign \U3/U5/DATA3_27  = NewElement[27];
  assign \U3/U5/DATA3_28  = NewElement[28];
  assign \U3/U5/DATA3_29  = NewElement[29];
  assign \U3/U5/DATA3_30  = NewElement[30];
  assign \U3/U5/DATA3_31  = NewElement[31];
  assign \U3/U5/DATA3_32  = NewElement[32];
  assign \U3/U5/DATA3_33  = NewElement[33];
  assign \U3/U5/DATA3_34  = NewElement[34];
  assign \U3/U5/DATA3_35  = NewElement[35];
  assign \U3/U5/DATA3_36  = NewElement[36];
  assign \U3/U5/DATA3_37  = NewElement[37];
  assign \U3/U5/DATA3_38  = NewElement[38];
  assign \U3/U5/DATA3_39  = NewElement[39];
  assign \U3/U5/DATA3_40  = NewElement[40];
  assign \U3/U5/DATA3_41  = NewElement[41];
  assign \U3/U5/DATA3_42  = NewElement[42];
  assign \U3/U5/DATA3_43  = NewElement[43];
  assign \U3/U5/DATA3_44  = NewElement[44];
  assign \U3/U5/DATA3_45  = NewElement[45];
  assign \U3/U5/DATA3_46  = NewElement[46];
  assign \U3/U5/DATA3_47  = NewElement[47];
  assign \U3/U5/DATA2_0  = NewDiagonalY[0];
  assign \U3/U5/DATA2_1  = NewDiagonalY[1];
  assign \U3/U5/DATA2_2  = NewDiagonalY[2];
  assign \U3/U5/DATA2_3  = NewDiagonalY[3];
  assign \U3/U5/DATA2_4  = NewDiagonalY[4];
  assign \U3/U5/DATA2_5  = NewDiagonalY[5];
  assign \U3/U5/DATA2_6  = NewDiagonalY[6];
  assign \U3/U5/DATA2_7  = NewDiagonalY[7];
  assign \U3/U5/DATA2_8  = NewDiagonalY[8];
  assign \U3/U5/DATA2_9  = NewDiagonalY[9];
  assign \U3/U5/DATA2_10  = NewDiagonalY[10];
  assign \U3/U5/DATA2_11  = NewDiagonalY[11];
  assign \U3/U5/DATA2_12  = NewDiagonalY[12];
  assign \U3/U5/DATA2_13  = NewDiagonalY[13];
  assign \U3/U5/DATA2_14  = NewDiagonalY[14];
  assign \U3/U5/DATA2_15  = NewDiagonalY[15];
  assign \U3/U5/DATA2_16  = NewDiagonalY[16];
  assign \U3/U5/DATA2_17  = NewDiagonalY[17];
  assign \U3/U5/DATA2_18  = NewDiagonalY[18];
  assign \U3/U5/DATA2_19  = NewDiagonalY[19];
  assign \U3/U5/DATA2_20  = NewDiagonalY[20];
  assign \U3/U5/DATA2_21  = NewDiagonalY[21];
  assign \U3/U5/DATA2_22  = NewDiagonalY[22];
  assign \U3/U5/DATA2_23  = NewDiagonalY[23];
  assign \U3/U5/DATA2_24  = NewDiagonalY[24];
  assign \U3/U5/DATA2_25  = NewDiagonalY[25];
  assign \U3/U5/DATA2_26  = NewDiagonalY[26];
  assign \U3/U5/DATA2_27  = NewDiagonalY[27];
  assign \U3/U5/DATA2_28  = NewDiagonalY[28];
  assign \U3/U5/DATA2_29  = NewDiagonalY[29];
  assign \U3/U5/DATA2_30  = NewDiagonalY[30];
  assign \U3/U5/DATA2_31  = NewDiagonalY[31];
  assign \U3/U5/DATA2_32  = NewDiagonalY[32];
  assign \U3/U5/DATA2_33  = NewDiagonalY[33];
  assign \U3/U5/DATA2_34  = NewDiagonalY[34];
  assign \U3/U5/DATA2_35  = NewDiagonalY[35];
  assign \U3/U5/DATA2_36  = NewDiagonalY[36];
  assign \U3/U5/DATA2_37  = NewDiagonalY[37];
  assign \U3/U5/DATA2_38  = NewDiagonalY[38];
  assign \U3/U5/DATA2_39  = NewDiagonalY[39];
  assign \U3/U5/DATA2_40  = NewDiagonalY[40];
  assign \U3/U5/DATA2_41  = NewDiagonalY[41];
  assign \U3/U5/DATA2_42  = NewDiagonalY[42];
  assign \U3/U5/DATA2_43  = NewDiagonalY[43];
  assign \U3/U5/DATA2_44  = NewDiagonalY[44];
  assign \U3/U5/DATA2_45  = NewDiagonalY[45];
  assign \U3/U5/DATA2_46  = NewDiagonalY[46];
  assign \U3/U5/DATA2_47  = NewDiagonalY[47];
  assign \U3/U5/DATA1_0  = NewDiagonalX[0];
  assign \U3/U5/DATA1_1  = NewDiagonalX[1];
  assign \U3/U5/DATA1_2  = NewDiagonalX[2];
  assign \U3/U5/DATA1_3  = NewDiagonalX[3];
  assign \U3/U5/DATA1_4  = NewDiagonalX[4];
  assign \U3/U5/DATA1_5  = NewDiagonalX[5];
  assign \U3/U5/DATA1_6  = NewDiagonalX[6];
  assign \U3/U5/DATA1_7  = NewDiagonalX[7];
  assign \U3/U5/DATA1_8  = NewDiagonalX[8];
  assign \U3/U5/DATA1_9  = NewDiagonalX[9];
  assign \U3/U5/DATA1_10  = NewDiagonalX[10];
  assign \U3/U5/DATA1_11  = NewDiagonalX[11];
  assign \U3/U5/DATA1_12  = NewDiagonalX[12];
  assign \U3/U5/DATA1_13  = NewDiagonalX[13];
  assign \U3/U5/DATA1_14  = NewDiagonalX[14];
  assign \U3/U5/DATA1_15  = NewDiagonalX[15];
  assign \U3/U5/DATA1_16  = NewDiagonalX[16];
  assign \U3/U5/DATA1_17  = NewDiagonalX[17];
  assign \U3/U5/DATA1_18  = NewDiagonalX[18];
  assign \U3/U5/DATA1_19  = NewDiagonalX[19];
  assign \U3/U5/DATA1_20  = NewDiagonalX[20];
  assign \U3/U5/DATA1_21  = NewDiagonalX[21];
  assign \U3/U5/DATA1_22  = NewDiagonalX[22];
  assign \U3/U5/DATA1_23  = NewDiagonalX[23];
  assign \U3/U5/DATA1_24  = NewDiagonalX[24];
  assign \U3/U5/DATA1_25  = NewDiagonalX[25];
  assign \U3/U5/DATA1_26  = NewDiagonalX[26];
  assign \U3/U5/DATA1_27  = NewDiagonalX[27];
  assign \U3/U5/DATA1_28  = NewDiagonalX[28];
  assign \U3/U5/DATA1_29  = NewDiagonalX[29];
  assign \U3/U5/DATA1_30  = NewDiagonalX[30];
  assign \U3/U5/DATA1_31  = NewDiagonalX[31];
  assign \U3/U5/DATA1_32  = NewDiagonalX[32];
  assign \U3/U5/DATA1_33  = NewDiagonalX[33];
  assign \U3/U5/DATA1_34  = NewDiagonalX[34];
  assign \U3/U5/DATA1_35  = NewDiagonalX[35];
  assign \U3/U5/DATA1_36  = NewDiagonalX[36];
  assign \U3/U5/DATA1_37  = NewDiagonalX[37];
  assign \U3/U5/DATA1_38  = NewDiagonalX[38];
  assign \U3/U5/DATA1_39  = NewDiagonalX[39];
  assign \U3/U5/DATA1_40  = NewDiagonalX[40];
  assign \U3/U5/DATA1_41  = NewDiagonalX[41];
  assign \U3/U5/DATA1_42  = NewDiagonalX[42];
  assign \U3/U5/DATA1_43  = NewDiagonalX[43];
  assign \U3/U5/DATA1_44  = NewDiagonalX[44];
  assign \U3/U5/DATA1_45  = NewDiagonalX[45];
  assign \U3/U5/DATA1_46  = NewDiagonalX[46];
  assign \U3/U5/DATA1_47  = NewDiagonalX[47];
  assign OutputReq1[0] = \U3/U7/Z_0 ;
  assign OutputReq1[1] = \U3/U7/Z_1 ;
  assign OutputReq1[2] = \U3/U7/Z_2 ;
  assign OutputReq1[3] = \U3/U7/Z_3 ;
  assign OutputReq1[4] = \U3/U7/Z_4 ;
  assign OutputReq1[5] = \U3/U7/Z_5 ;
  assign OutputReq1[6] = \U3/U7/Z_6 ;
  assign OutputReq1[7] = \U3/U7/Z_7 ;
  assign OutputReq1[8] = \U3/U7/Z_8 ;
  assign OutputReq1[9] = \U3/U7/Z_9 ;
  assign OutputReq1[10] = \U3/U7/Z_10 ;
  assign \U3/U7/DATA7_0  = ComputeReq[0];
  assign \U3/U7/DATA7_1  = ComputeReq[1];
  assign \U3/U7/DATA7_2  = ComputeReq[2];
  assign \U3/U7/DATA7_3  = ComputeReq[3];
  assign \U3/U7/DATA7_4  = ComputeReq[4];
  assign \U3/U7/DATA7_5  = ComputeReq[5];
  assign \U3/U7/DATA7_6  = ComputeReq[6];
  assign \U3/U7/DATA7_7  = ComputeReq[7];
  assign \U3/U7/DATA7_8  = ComputeReq[8];
  assign \U3/U7/DATA7_9  = ComputeReq[9];
  assign \U3/U7/DATA7_10  = ComputeReq[10];
  assign \U3/U7/DATA6_0  = PosRowY[2];
  assign \U3/U7/DATA6_1  = PosRowY[3];
  assign \U3/U7/DATA6_2  = PosRowY[4];
  assign \U3/U7/DATA6_3  = PosRowY[5];
  assign \U3/U7/DATA6_4  = PosRowY[6];
  assign \U3/U7/DATA6_5  = PosRowY[7];
  assign \U3/U7/DATA6_6  = PosRowY[8];
  assign \U3/U7/DATA6_7  = PosRowY[9];
  assign \U3/U7/DATA6_8  = PosRowY[10];
  assign \U3/U7/DATA6_9  = PosRowY[11];
  assign \U3/U7/DATA6_10  = PosRowY[12];
  assign \U3/U7/DATA5_0  = PosRowX[2];
  assign \U3/U7/DATA5_1  = PosRowX[3];
  assign \U3/U7/DATA5_2  = PosRowX[4];
  assign \U3/U7/DATA5_3  = PosRowX[5];
  assign \U3/U7/DATA5_4  = PosRowX[6];
  assign \U3/U7/DATA5_5  = PosRowX[7];
  assign \U3/U7/DATA5_6  = PosRowX[8];
  assign \U3/U7/DATA5_7  = PosRowX[9];
  assign \U3/U7/DATA5_8  = PosRowX[10];
  assign \U3/U7/DATA5_9  = PosRowX[11];
  assign \U3/U7/DATA5_10  = PosRowX[12];
  assign \U3/U7/DATA4_0  = PosDY[2];
  assign \U3/U7/DATA4_1  = PosDY[3];
  assign \U3/U7/DATA4_2  = PosDY[4];
  assign \U3/U7/DATA4_3  = PosDY[5];
  assign \U3/U7/DATA4_4  = PosDY[6];
  assign \U3/U7/DATA4_5  = PosDY[7];
  assign \U3/U7/DATA4_6  = PosDY[8];
  assign \U3/U7/DATA4_7  = PosDY[9];
  assign \U3/U7/DATA4_8  = PosDY[10];
  assign \U3/U7/DATA4_9  = PosDY[11];
  assign \U3/U7/DATA4_10  = PosDY[12];
  assign \U3/U7/DATA3_0  = PosDX[2];
  assign \U3/U7/DATA3_1  = PosDX[3];
  assign \U3/U7/DATA3_2  = PosDX[4];
  assign \U3/U7/DATA3_3  = PosDX[5];
  assign \U3/U7/DATA3_4  = PosDX[6];
  assign \U3/U7/DATA3_5  = PosDX[7];
  assign \U3/U7/DATA3_6  = PosDX[8];
  assign \U3/U7/DATA3_7  = PosDX[9];
  assign \U3/U7/DATA3_8  = PosDX[10];
  assign \U3/U7/DATA3_9  = PosDX[11];
  assign \U3/U7/DATA3_10  = PosDX[12];
  assign \U3/U7/DATA2_0  = Update_2Req1[0];
  assign \U3/U7/DATA2_1  = Update_2Req1[1];
  assign \U3/U7/DATA2_2  = Update_2Req1[2];
  assign \U3/U7/DATA2_3  = Update_2Req1[3];
  assign \U3/U7/DATA2_4  = Update_2Req1[4];
  assign \U3/U7/DATA2_5  = Update_2Req1[5];
  assign \U3/U7/DATA2_6  = Update_2Req1[6];
  assign \U3/U7/DATA2_7  = Update_2Req1[7];
  assign \U3/U7/DATA2_8  = Update_2Req1[8];
  assign \U3/U7/DATA2_9  = Update_2Req1[9];
  assign \U3/U7/DATA2_10  = Update_2Req1[10];
  assign \U3/U7/DATA1_0  = Update_1Req1[0];
  assign \U3/U7/DATA1_1  = Update_1Req1[1];
  assign \U3/U7/DATA1_2  = Update_1Req1[2];
  assign \U3/U7/DATA1_3  = Update_1Req1[3];
  assign \U3/U7/DATA1_4  = Update_1Req1[4];
  assign \U3/U7/DATA1_5  = Update_1Req1[5];
  assign \U3/U7/DATA1_6  = Update_1Req1[6];
  assign \U3/U7/DATA1_7  = Update_1Req1[7];
  assign \U3/U7/DATA1_8  = Update_1Req1[8];
  assign \U3/U7/DATA1_9  = Update_1Req1[9];
  assign \U3/U7/DATA1_10  = Update_1Req1[10];
  assign ArbiterPos[0] = \U3/U8/Z_0 ;
  assign ArbiterPos[1] = \U3/U8/Z_1 ;
  assign \U3/U8/DATA4_0  = PosRowY[0];
  assign \U3/U8/DATA4_1  = PosRowY[1];
  assign \U3/U8/DATA3_0  = PosRowX[0];
  assign \U3/U8/DATA3_1  = PosRowX[1];
  assign \U3/U8/DATA2_0  = PosDY[0];
  assign \U3/U8/DATA2_1  = PosDY[1];
  assign \U3/U8/DATA1_0  = PosDX[0];
  assign \U3/U8/DATA1_1  = PosDX[1];
  assign WriteReq[0] = \U3/U9/Z_0 ;
  assign WriteReq[1] = \U3/U9/Z_1 ;
  assign WriteReq[2] = \U3/U9/Z_2 ;
  assign WriteReq[3] = \U3/U9/Z_3 ;
  assign WriteReq[4] = \U3/U9/Z_4 ;
  assign WriteReq[5] = \U3/U9/Z_5 ;
  assign WriteReq[6] = \U3/U9/Z_6 ;
  assign WriteReq[7] = \U3/U9/Z_7 ;
  assign WriteReq[8] = \U3/U9/Z_8 ;
  assign WriteReq[9] = \U3/U9/Z_9 ;
  assign WriteReq[10] = \U3/U9/Z_10 ;
  assign \U3/U10/DATA3_0  = DiagonalDoneX;
  assign \U3/U10/DATA1_0  = EnableChange;

  DFF_X1 \current_state_reg[1]  ( .D(\U4/Z_1 ), .CK(clock), .Q(n1828), .QN(n8)
         );
  NAND3_X2 U5 ( .A1(n4801), .A2(n39), .A3(n4770), .ZN(n38) );
  NOR2_X2 U7 ( .A1(n4770), .A2(n42), .ZN(n41) );
  OAI22_X2 U8 ( .A1(reset), .A2(n43), .B1(n44), .B2(n2961), .ZN(\U4/Z_1 ) );
  NOR2_X2 U9 ( .A1(n1830), .A2(reset), .ZN(n39) );
  NOR3_X2 U11 ( .A1(n4800), .A2(n4770), .A3(\U3/U4/DATA2_0 ), .ZN(n46) );
  NOR2_X2 U12 ( .A1(n4771), .A2(reset), .ZN(\U4/Z_0 ) );
  NAND3_X2 U14 ( .A1(n50), .A2(n4768), .A3(n1830), .ZN(n37) );
  NAND3_X2 U16 ( .A1(n4799), .A2(n4768), .A3(\U3/U10/DATA1_0 ), .ZN(n49) );
  AOI221_X2 U17 ( .B1(\U3/U10/DATA3_0 ), .B2(n4798), .C1(n4770), .C2(n52), .A(
        n53), .ZN(n48) );
  NOR3_X2 U18 ( .A1(n42), .A2(n4770), .A3(\U3/U4/DATA2_0 ), .ZN(n53) );
  OAI221_X2 U19 ( .B1(n2960), .B2(n54), .C1(n55), .C2(n45), .A(n56), .ZN(n52)
         );
  NAND2_X2 U20 ( .A1(n57), .A2(n58), .ZN(n45) );
  NOR4_X2 U21 ( .A1(n59), .A2(\U3/U7/DATA6_5 ), .A3(\U3/U7/DATA6_7 ), .A4(
        \U3/U7/DATA6_6 ), .ZN(n58) );
  NOR4_X2 U22 ( .A1(n60), .A2(\U3/U7/DATA6_0 ), .A3(\U3/U7/DATA6_10 ), .A4(
        \U3/U7/DATA6_1 ), .ZN(n57) );
  NOR3_X2 U23 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n54) );
  OAI221_X2 U24 ( .B1(n51), .B2(n4790), .C1(n4770), .C2(n4779), .A(n65), .ZN(
        \U3/U9/Z_7 ) );
  OAI221_X2 U26 ( .B1(n51), .B2(n4791), .C1(n4770), .C2(n4780), .A(n66), .ZN(
        \U3/U9/Z_6 ) );
  OAI221_X2 U28 ( .B1(n51), .B2(n4792), .C1(n4770), .C2(n4781), .A(n67), .ZN(
        \U3/U9/Z_5 ) );
  OAI221_X2 U30 ( .B1(n51), .B2(n4793), .C1(n4770), .C2(n4782), .A(n68), .ZN(
        \U3/U9/Z_4 ) );
  OAI221_X2 U32 ( .B1(n51), .B2(n4794), .C1(n4770), .C2(n4783), .A(n69), .ZN(
        \U3/U9/Z_3 ) );
  OAI221_X2 U34 ( .B1(n51), .B2(n4795), .C1(n4770), .C2(n4784), .A(n70), .ZN(
        \U3/U9/Z_2 ) );
  OAI221_X2 U36 ( .B1(n51), .B2(n4796), .C1(n4770), .C2(n4785), .A(n71), .ZN(
        \U3/U9/Z_1 ) );
  OAI221_X2 U38 ( .B1(n51), .B2(n4797), .C1(n4770), .C2(n4786), .A(n72), .ZN(
        \U3/U9/Z_0 ) );
  OAI221_X2 U40 ( .B1(n51), .B2(n4787), .C1(n4770), .C2(n4776), .A(n73), .ZN(
        \U3/U9/Z_10 ) );
  OAI221_X2 U42 ( .B1(n51), .B2(n4788), .C1(n4770), .C2(n4777), .A(n74), .ZN(
        \U3/U9/Z_9 ) );
  OAI221_X2 U44 ( .B1(n51), .B2(n4789), .C1(n4770), .C2(n4778), .A(n75), .ZN(
        \U3/U9/Z_8 ) );
  OAI221_X2 U46 ( .B1(n56), .B2(n4772), .C1(n55), .C2(n4774), .A(n76), .ZN(
        \U3/U8/Z_1 ) );
  OAI221_X2 U48 ( .B1(n56), .B2(n4773), .C1(n55), .C2(n4775), .A(n77), .ZN(
        \U3/U8/Z_0 ) );
  NAND3_X2 U50 ( .A1(n78), .A2(n79), .A3(n80), .ZN(\U3/U7/Z_9 ) );
  NAND3_X2 U54 ( .A1(n86), .A2(n87), .A3(n88), .ZN(\U3/U7/Z_8 ) );
  NAND3_X2 U58 ( .A1(n89), .A2(n90), .A3(n91), .ZN(\U3/U7/Z_7 ) );
  NAND3_X2 U62 ( .A1(n92), .A2(n93), .A3(n94), .ZN(\U3/U7/Z_6 ) );
  NAND3_X2 U66 ( .A1(n95), .A2(n96), .A3(n97), .ZN(\U3/U7/Z_5 ) );
  NAND3_X2 U70 ( .A1(n98), .A2(n99), .A3(n100), .ZN(\U3/U7/Z_4 ) );
  NAND3_X2 U74 ( .A1(n101), .A2(n102), .A3(n103), .ZN(\U3/U7/Z_3 ) );
  NAND3_X2 U78 ( .A1(n104), .A2(n105), .A3(n106), .ZN(\U3/U7/Z_2 ) );
  NAND3_X2 U82 ( .A1(n107), .A2(n108), .A3(n109), .ZN(\U3/U7/Z_10 ) );
  NAND3_X2 U86 ( .A1(n110), .A2(n111), .A3(n112), .ZN(\U3/U7/Z_1 ) );
  NAND3_X2 U90 ( .A1(n113), .A2(n114), .A3(n115), .ZN(\U3/U7/Z_0 ) );
  INV_X4 U98 ( .A(n116), .ZN(\U3/U5/Z_9 ) );
  INV_X4 U100 ( .A(n118), .ZN(\U3/U5/Z_8 ) );
  INV_X4 U102 ( .A(n119), .ZN(\U3/U5/Z_7 ) );
  INV_X4 U104 ( .A(n120), .ZN(\U3/U5/Z_6 ) );
  INV_X4 U106 ( .A(n121), .ZN(\U3/U5/Z_5 ) );
  INV_X4 U108 ( .A(n122), .ZN(\U3/U5/Z_47 ) );
  INV_X4 U110 ( .A(n123), .ZN(\U3/U5/Z_46 ) );
  INV_X4 U112 ( .A(n124), .ZN(\U3/U5/Z_45 ) );
  INV_X4 U114 ( .A(n125), .ZN(\U3/U5/Z_44 ) );
  INV_X4 U116 ( .A(n126), .ZN(\U3/U5/Z_43 ) );
  INV_X4 U118 ( .A(n127), .ZN(\U3/U5/Z_42 ) );
  INV_X4 U120 ( .A(n128), .ZN(\U3/U5/Z_41 ) );
  INV_X4 U122 ( .A(n129), .ZN(\U3/U5/Z_40 ) );
  INV_X4 U124 ( .A(n130), .ZN(\U3/U5/Z_4 ) );
  INV_X4 U126 ( .A(n131), .ZN(\U3/U5/Z_39 ) );
  INV_X4 U128 ( .A(n132), .ZN(\U3/U5/Z_38 ) );
  INV_X4 U130 ( .A(n133), .ZN(\U3/U5/Z_37 ) );
  INV_X4 U132 ( .A(n134), .ZN(\U3/U5/Z_36 ) );
  INV_X4 U134 ( .A(n135), .ZN(\U3/U5/Z_35 ) );
  INV_X4 U136 ( .A(n136), .ZN(\U3/U5/Z_34 ) );
  INV_X4 U138 ( .A(n137), .ZN(\U3/U5/Z_33 ) );
  INV_X4 U140 ( .A(n138), .ZN(\U3/U5/Z_32 ) );
  INV_X4 U142 ( .A(n139), .ZN(\U3/U5/Z_31 ) );
  INV_X4 U144 ( .A(n140), .ZN(\U3/U5/Z_30 ) );
  INV_X4 U146 ( .A(n141), .ZN(\U3/U5/Z_3 ) );
  INV_X4 U148 ( .A(n142), .ZN(\U3/U5/Z_29 ) );
  INV_X4 U150 ( .A(n143), .ZN(\U3/U5/Z_28 ) );
  INV_X4 U152 ( .A(n144), .ZN(\U3/U5/Z_27 ) );
  INV_X4 U154 ( .A(n145), .ZN(\U3/U5/Z_26 ) );
  INV_X4 U156 ( .A(n146), .ZN(\U3/U5/Z_25 ) );
  INV_X4 U158 ( .A(n147), .ZN(\U3/U5/Z_24 ) );
  INV_X4 U160 ( .A(n148), .ZN(\U3/U5/Z_23 ) );
  INV_X4 U162 ( .A(n149), .ZN(\U3/U5/Z_22 ) );
  INV_X4 U164 ( .A(n150), .ZN(\U3/U5/Z_21 ) );
  INV_X4 U166 ( .A(n151), .ZN(\U3/U5/Z_20 ) );
  INV_X4 U168 ( .A(n152), .ZN(\U3/U5/Z_2 ) );
  INV_X4 U170 ( .A(n153), .ZN(\U3/U5/Z_19 ) );
  INV_X4 U172 ( .A(n154), .ZN(\U3/U5/Z_18 ) );
  INV_X4 U174 ( .A(n155), .ZN(\U3/U5/Z_17 ) );
  INV_X4 U176 ( .A(n156), .ZN(\U3/U5/Z_16 ) );
  INV_X4 U178 ( .A(n157), .ZN(\U3/U5/Z_15 ) );
  INV_X4 U180 ( .A(n158), .ZN(\U3/U5/Z_14 ) );
  INV_X4 U182 ( .A(n159), .ZN(\U3/U5/Z_13 ) );
  INV_X4 U184 ( .A(n160), .ZN(\U3/U5/Z_12 ) );
  INV_X4 U186 ( .A(n161), .ZN(\U3/U5/Z_11 ) );
  INV_X4 U188 ( .A(n162), .ZN(\U3/U5/Z_10 ) );
  INV_X4 U190 ( .A(n163), .ZN(\U3/U5/Z_1 ) );
  INV_X4 U192 ( .A(n164), .ZN(\U3/U5/Z_0 ) );
  NAND2_X2 U195 ( .A1(n1828), .A2(n4800), .ZN(n56) );
  NAND2_X2 U196 ( .A1(n2960), .A2(n8), .ZN(n55) );
  INV_X4 U198 ( .A(n165), .ZN(\U3/U3/Z_9 ) );
  INV_X4 U200 ( .A(n166), .ZN(\U3/U3/Z_8 ) );
  INV_X4 U202 ( .A(n167), .ZN(\U3/U3/Z_7 ) );
  INV_X4 U204 ( .A(n168), .ZN(\U3/U3/Z_6 ) );
  INV_X4 U206 ( .A(n169), .ZN(\U3/U3/Z_5 ) );
  INV_X4 U208 ( .A(n170), .ZN(\U3/U3/Z_4 ) );
  INV_X4 U210 ( .A(n171), .ZN(\U3/U3/Z_3 ) );
  INV_X4 U212 ( .A(n172), .ZN(\U3/U3/Z_2 ) );
  INV_X4 U214 ( .A(n173), .ZN(\U3/U3/Z_10 ) );
  INV_X4 U216 ( .A(n174), .ZN(\U3/U3/Z_1 ) );
  INV_X4 U218 ( .A(n175), .ZN(\U3/U3/Z_0 ) );
  INV_X4 U220 ( .A(n43), .ZN(\U3/U2/Z_0 ) );
  NAND2_X2 U221 ( .A1(n82), .A2(n2960), .ZN(n43) );
  NAND2_X2 U224 ( .A1(n1828), .A2(n2960), .ZN(n42) );
  OR4_X1 U258 ( .A1(\U3/U7/DATA6_8 ), .A2(\U3/U7/DATA6_9 ), .A3(
        \U3/U8/DATA4_0 ), .A4(\U3/U8/DATA4_1 ), .ZN(n59) );
  OR3_X1 U259 ( .A1(\U3/U7/DATA6_3 ), .A2(\U3/U7/DATA6_4 ), .A3(
        \U3/U7/DATA6_2 ), .ZN(n60) );
  OR3_X1 U260 ( .A1(\U3/U7/DATA5_6 ), .A2(\U3/U7/DATA5_7 ), .A3(
        \U3/U7/DATA5_5 ), .ZN(n63) );
  OR4_X1 U261 ( .A1(\U3/U7/DATA5_8 ), .A2(\U3/U7/DATA5_9 ), .A3(
        \U3/U8/DATA3_0 ), .A4(\U3/U8/DATA3_1 ), .ZN(n62) );
  OR4_X1 U262 ( .A1(\U3/U7/DATA5_1 ), .A2(\U3/U7/DATA5_10 ), .A3(
        \U3/U7/DATA5_0 ), .A4(n64), .ZN(n61) );
  OR3_X1 U263 ( .A1(\U3/U7/DATA5_2 ), .A2(\U3/U7/DATA5_4 ), .A3(
        \U3/U7/DATA5_3 ), .ZN(n64) );
  DFF_X2 \current_state_reg[3]  ( .D(\U4/Z_3 ), .CK(clock), .Q(n1830) );
  DFF_X2 \current_state_reg[2]  ( .D(n2962), .CK(clock), .Q(n4770), .QN(n2959)
         );
  DFF_X2 \current_state_reg[0]  ( .D(\U4/Z_0 ), .CK(clock), .Q(n2960), .QN(
        CompStart) );
  NAND2_X4 U3 ( .A1(n55), .A2(n56), .ZN(n2958) );
  NOR2_X1 U4 ( .A1(n40), .A2(n2961), .ZN(n2962) );
  INV_X1 U6 ( .A(n39), .ZN(n2961) );
  BUF_X4 U10 ( .A(Row1[11]), .Z(Output_1Row1[11]) );
  BUF_X4 U13 ( .A(Row1[12]), .Z(Output_1Row1[12]) );
  BUF_X4 U15 ( .A(Row1[13]), .Z(Output_1Row1[13]) );
  BUF_X4 U25 ( .A(Row1[14]), .Z(Output_1Row1[14]) );
  BUF_X4 U27 ( .A(Row1[15]), .Z(Output_1Row1[15]) );
  BUF_X4 U29 ( .A(Row1[27]), .Z(Output_1Row1[27]) );
  BUF_X4 U31 ( .A(Row1[28]), .Z(Output_1Row1[28]) );
  BUF_X4 U33 ( .A(Row1[29]), .Z(Output_1Row1[29]) );
  BUF_X4 U35 ( .A(Row1[30]), .Z(Output_1Row1[30]) );
  BUF_X4 U37 ( .A(Row1[31]), .Z(Output_1Row1[31]) );
  BUF_X4 U39 ( .A(Row1[43]), .Z(Output_1Row1[43]) );
  BUF_X4 U41 ( .A(Row1[44]), .Z(Output_1Row1[44]) );
  BUF_X4 U43 ( .A(Row1[45]), .Z(Output_1Row1[45]) );
  BUF_X4 U45 ( .A(Row1[46]), .Z(Output_1Row1[46]) );
  BUF_X4 U47 ( .A(Row1[47]), .Z(Output_1Row1[47]) );
  BUF_X4 U49 ( .A(Row1[75]), .Z(Output_1Row1[75]) );
  BUF_X4 U51 ( .A(Row1[76]), .Z(Output_1Row1[76]) );
  BUF_X4 U52 ( .A(Row1[77]), .Z(Output_1Row1[77]) );
  BUF_X4 U53 ( .A(Row1[78]), .Z(Output_1Row1[78]) );
  BUF_X4 U55 ( .A(Row1[79]), .Z(Output_1Row1[79]) );
  BUF_X4 U56 ( .A(Row1[91]), .Z(Output_1Row1[91]) );
  BUF_X4 U57 ( .A(Row1[92]), .Z(Output_1Row1[92]) );
  BUF_X4 U59 ( .A(Row1[93]), .Z(Output_1Row1[93]) );
  BUF_X4 U60 ( .A(Row1[94]), .Z(Output_1Row1[94]) );
  BUF_X4 U61 ( .A(Row1[95]), .Z(Output_1Row1[95]) );
  BUF_X4 U63 ( .A(Row1[107]), .Z(Output_1Row1[107]) );
  BUF_X4 U64 ( .A(Row1[108]), .Z(Output_1Row1[108]) );
  BUF_X4 U65 ( .A(Row1[109]), .Z(Output_1Row1[109]) );
  BUF_X4 U67 ( .A(Row1[110]), .Z(Output_1Row1[110]) );
  BUF_X4 U68 ( .A(Row1[111]), .Z(Output_1Row1[111]) );
  BUF_X4 U69 ( .A(Row1[139]), .Z(Output_1Row1[139]) );
  BUF_X4 U71 ( .A(Row1[140]), .Z(Output_1Row1[140]) );
  BUF_X4 U72 ( .A(Row1[141]), .Z(Output_1Row1[141]) );
  BUF_X4 U73 ( .A(Row1[142]), .Z(Output_1Row1[142]) );
  BUF_X4 U75 ( .A(Row1[143]), .Z(Output_1Row1[143]) );
  BUF_X4 U76 ( .A(Row1[155]), .Z(Output_1Row1[155]) );
  BUF_X4 U77 ( .A(Row1[156]), .Z(Output_1Row1[156]) );
  BUF_X4 U79 ( .A(Row1[157]), .Z(Output_1Row1[157]) );
  BUF_X4 U80 ( .A(Row1[158]), .Z(Output_1Row1[158]) );
  BUF_X4 U81 ( .A(Row1[159]), .Z(Output_1Row1[159]) );
  BUF_X4 U83 ( .A(Row1[171]), .Z(Output_1Row1[171]) );
  BUF_X4 U84 ( .A(Row1[172]), .Z(Output_1Row1[172]) );
  BUF_X4 U85 ( .A(Row1[173]), .Z(Output_1Row1[173]) );
  BUF_X4 U87 ( .A(Row1[174]), .Z(Output_1Row1[174]) );
  BUF_X4 U88 ( .A(Row1[175]), .Z(Output_1Row1[175]) );
  BUF_X4 U89 ( .A(Row1[203]), .Z(Output_1Row1[203]) );
  BUF_X4 U91 ( .A(Row1[204]), .Z(Output_1Row1[204]) );
  BUF_X4 U92 ( .A(Row1[205]), .Z(Output_1Row1[205]) );
  BUF_X4 U93 ( .A(Row1[206]), .Z(Output_1Row1[206]) );
  BUF_X4 U94 ( .A(Row1[207]), .Z(Output_1Row1[207]) );
  BUF_X4 U95 ( .A(Row1[219]), .Z(Output_1Row1[219]) );
  BUF_X4 U96 ( .A(Row1[220]), .Z(Output_1Row1[220]) );
  BUF_X4 U97 ( .A(Row1[221]), .Z(Output_1Row1[221]) );
  BUF_X4 U99 ( .A(Row1[222]), .Z(Output_1Row1[222]) );
  BUF_X4 U101 ( .A(Row1[223]), .Z(Output_1Row1[223]) );
  BUF_X4 U103 ( .A(Row1[235]), .Z(Output_1Row1[235]) );
  BUF_X4 U105 ( .A(Row1[236]), .Z(Output_1Row1[236]) );
  BUF_X4 U107 ( .A(Row1[237]), .Z(Output_1Row1[237]) );
  BUF_X4 U109 ( .A(Row1[238]), .Z(Output_1Row1[238]) );
  BUF_X4 U111 ( .A(Row1[239]), .Z(Output_1Row1[239]) );
  BUF_X4 U113 ( .A(Row2[11]), .Z(Output_1Row2[11]) );
  BUF_X4 U115 ( .A(Row2[12]), .Z(Output_1Row2[12]) );
  BUF_X4 U117 ( .A(Row2[13]), .Z(Output_1Row2[13]) );
  BUF_X4 U119 ( .A(Row2[14]), .Z(Output_1Row2[14]) );
  BUF_X4 U121 ( .A(Row2[15]), .Z(Output_1Row2[15]) );
  BUF_X4 U123 ( .A(Row2[27]), .Z(Output_1Row2[27]) );
  BUF_X4 U125 ( .A(Row2[28]), .Z(Output_1Row2[28]) );
  BUF_X4 U127 ( .A(Row2[29]), .Z(Output_1Row2[29]) );
  BUF_X4 U129 ( .A(Row2[30]), .Z(Output_1Row2[30]) );
  BUF_X4 U131 ( .A(Row2[31]), .Z(Output_1Row2[31]) );
  BUF_X4 U133 ( .A(Row2[43]), .Z(Output_1Row2[43]) );
  BUF_X4 U135 ( .A(Row2[44]), .Z(Output_1Row2[44]) );
  BUF_X4 U137 ( .A(Row2[45]), .Z(Output_1Row2[45]) );
  BUF_X4 U139 ( .A(Row2[46]), .Z(Output_1Row2[46]) );
  BUF_X4 U141 ( .A(Row2[47]), .Z(Output_1Row2[47]) );
  BUF_X4 U143 ( .A(Row2[59]), .Z(Output_1Row2[59]) );
  BUF_X4 U145 ( .A(Row2[60]), .Z(Output_1Row2[60]) );
  BUF_X4 U147 ( .A(Row2[61]), .Z(Output_1Row2[61]) );
  BUF_X4 U149 ( .A(Row2[62]), .Z(Output_1Row2[62]) );
  BUF_X4 U151 ( .A(Row2[63]), .Z(Output_1Row2[63]) );
  BUF_X4 U153 ( .A(Row2[75]), .Z(Output_1Row2[75]) );
  BUF_X4 U155 ( .A(Row2[76]), .Z(Output_1Row2[76]) );
  BUF_X4 U157 ( .A(Row2[77]), .Z(Output_1Row2[77]) );
  BUF_X4 U159 ( .A(Row2[78]), .Z(Output_1Row2[78]) );
  BUF_X4 U161 ( .A(Row2[79]), .Z(Output_1Row2[79]) );
  BUF_X4 U163 ( .A(Row2[91]), .Z(Output_1Row2[91]) );
  BUF_X4 U165 ( .A(Row2[92]), .Z(Output_1Row2[92]) );
  BUF_X4 U167 ( .A(Row2[93]), .Z(Output_1Row2[93]) );
  BUF_X4 U169 ( .A(Row2[94]), .Z(Output_1Row2[94]) );
  BUF_X4 U171 ( .A(Row2[95]), .Z(Output_1Row2[95]) );
  BUF_X4 U173 ( .A(Row2[107]), .Z(Output_1Row2[107]) );
  BUF_X4 U175 ( .A(Row2[108]), .Z(Output_1Row2[108]) );
  BUF_X4 U177 ( .A(Row2[109]), .Z(Output_1Row2[109]) );
  BUF_X4 U179 ( .A(Row2[110]), .Z(Output_1Row2[110]) );
  BUF_X4 U181 ( .A(Row2[111]), .Z(Output_1Row2[111]) );
  BUF_X4 U183 ( .A(Row2[123]), .Z(Output_1Row2[123]) );
  BUF_X4 U185 ( .A(Row2[124]), .Z(Output_1Row2[124]) );
  BUF_X4 U187 ( .A(Row2[125]), .Z(Output_1Row2[125]) );
  BUF_X4 U189 ( .A(Row2[126]), .Z(Output_1Row2[126]) );
  BUF_X4 U191 ( .A(Row2[127]), .Z(Output_1Row2[127]) );
  BUF_X4 U193 ( .A(Row2[139]), .Z(Output_1Row2[139]) );
  BUF_X4 U194 ( .A(Row2[140]), .Z(Output_1Row2[140]) );
  BUF_X4 U197 ( .A(Row2[141]), .Z(Output_1Row2[141]) );
  BUF_X4 U199 ( .A(Row2[142]), .Z(Output_1Row2[142]) );
  BUF_X4 U201 ( .A(Row2[143]), .Z(Output_1Row2[143]) );
  BUF_X4 U203 ( .A(Row2[155]), .Z(Output_1Row2[155]) );
  BUF_X4 U205 ( .A(Row2[156]), .Z(Output_1Row2[156]) );
  BUF_X4 U207 ( .A(Row2[157]), .Z(Output_1Row2[157]) );
  BUF_X4 U209 ( .A(Row2[158]), .Z(Output_1Row2[158]) );
  BUF_X4 U211 ( .A(Row2[159]), .Z(Output_1Row2[159]) );
  BUF_X4 U213 ( .A(Row2[171]), .Z(Output_1Row2[171]) );
  BUF_X4 U215 ( .A(Row2[172]), .Z(Output_1Row2[172]) );
  BUF_X4 U217 ( .A(Row2[173]), .Z(Output_1Row2[173]) );
  BUF_X4 U219 ( .A(Row2[174]), .Z(Output_1Row2[174]) );
  BUF_X4 U222 ( .A(Row2[175]), .Z(Output_1Row2[175]) );
  BUF_X4 U223 ( .A(Row2[187]), .Z(Output_1Row2[187]) );
  BUF_X4 U225 ( .A(Row2[188]), .Z(Output_1Row2[188]) );
  BUF_X4 U226 ( .A(Row2[189]), .Z(Output_1Row2[189]) );
  BUF_X4 U227 ( .A(Row2[190]), .Z(Output_1Row2[190]) );
  BUF_X4 U228 ( .A(Row2[191]), .Z(Output_1Row2[191]) );
  BUF_X4 U229 ( .A(Row2[203]), .Z(Output_1Row2[203]) );
  BUF_X4 U230 ( .A(Row2[204]), .Z(Output_1Row2[204]) );
  BUF_X4 U231 ( .A(Row2[205]), .Z(Output_1Row2[205]) );
  BUF_X4 U232 ( .A(Row2[206]), .Z(Output_1Row2[206]) );
  BUF_X4 U233 ( .A(Row2[207]), .Z(Output_1Row2[207]) );
  BUF_X4 U234 ( .A(Row2[219]), .Z(Output_1Row2[219]) );
  BUF_X4 U235 ( .A(Row2[220]), .Z(Output_1Row2[220]) );
  BUF_X4 U236 ( .A(Row2[221]), .Z(Output_1Row2[221]) );
  BUF_X4 U237 ( .A(Row2[222]), .Z(Output_1Row2[222]) );
  BUF_X4 U238 ( .A(Row2[223]), .Z(Output_1Row2[223]) );
  BUF_X4 U239 ( .A(Row2[235]), .Z(Output_1Row2[235]) );
  BUF_X4 U240 ( .A(Row2[236]), .Z(Output_1Row2[236]) );
  BUF_X4 U241 ( .A(Row2[237]), .Z(Output_1Row2[237]) );
  BUF_X4 U242 ( .A(Row2[238]), .Z(Output_1Row2[238]) );
  BUF_X4 U243 ( .A(Row2[239]), .Z(Output_1Row2[239]) );
  BUF_X4 U244 ( .A(Row2[251]), .Z(Output_1Row2[251]) );
  BUF_X4 U245 ( .A(Row2[252]), .Z(Output_1Row2[252]) );
  BUF_X4 U246 ( .A(Row2[253]), .Z(Output_1Row2[253]) );
  BUF_X4 U247 ( .A(Row2[254]), .Z(Output_1Row2[254]) );
  BUF_X4 U248 ( .A(Row2[255]), .Z(Output_1Row2[255]) );
  INV_X4 U249 ( .A(n4770), .ZN(n4768) );
  NOR2_X2 U250 ( .A1(n4768), .A2(n4800), .ZN(n84) );
  BUF_X4 U251 ( .A(Row1[54]), .Z(Output_2Row1[54]) );
  BUF_X4 U252 ( .A(Row1[55]), .Z(Output_2Row1[55]) );
  BUF_X4 U253 ( .A(Row1[118]), .Z(Output_2Row1[118]) );
  BUF_X4 U254 ( .A(Row1[119]), .Z(Output_2Row1[119]) );
  BUF_X4 U255 ( .A(Row1[50]), .Z(Output_2Row1[50]) );
  BUF_X4 U256 ( .A(Row1[49]), .Z(Output_2Row1[49]) );
  BUF_X4 U257 ( .A(Row1[51]), .Z(Output_2Row1[51]) );
  BUF_X4 U264 ( .A(Row1[53]), .Z(Output_2Row1[53]) );
  BUF_X4 U265 ( .A(Row1[115]), .Z(Output_2Row1[115]) );
  BUF_X4 U266 ( .A(Row1[114]), .Z(Output_2Row1[114]) );
  BUF_X4 U267 ( .A(Row1[62]), .Z(Output_2Row1[62]) );
  BUF_X4 U268 ( .A(Row1[126]), .Z(Output_2Row1[126]) );
  BUF_X4 U269 ( .A(Row1[61]), .Z(Output_2Row1[61]) );
  BUF_X4 U270 ( .A(Row1[63]), .Z(Output_2Row1[63]) );
  BUF_X4 U271 ( .A(Row1[127]), .Z(Output_2Row1[127]) );
  BUF_X4 U272 ( .A(Row1[182]), .Z(Output_2Row1[182]) );
  BUF_X4 U273 ( .A(Row1[183]), .Z(Output_2Row1[183]) );
  BUF_X4 U274 ( .A(Row1[48]), .Z(Output_2Row1[48]) );
  BUF_X4 U275 ( .A(Row1[52]), .Z(Output_2Row1[52]) );
  BUF_X4 U276 ( .A(Row1[178]), .Z(Output_2Row1[178]) );
  BUF_X4 U277 ( .A(Row1[181]), .Z(Output_2Row1[181]) );
  BUF_X4 U278 ( .A(Row1[180]), .Z(Output_2Row1[180]) );
  BUF_X4 U279 ( .A(Row1[112]), .Z(Output_2Row1[112]) );
  BUF_X4 U280 ( .A(Row1[117]), .Z(Output_2Row1[117]) );
  BUF_X4 U281 ( .A(Row1[116]), .Z(Output_2Row1[116]) );
  BUF_X4 U282 ( .A(Row1[179]), .Z(Output_2Row1[179]) );
  BUF_X4 U283 ( .A(Row1[177]), .Z(Output_2Row1[177]) );
  BUF_X4 U284 ( .A(Row1[176]), .Z(Output_2Row1[176]) );
  BUF_X4 U285 ( .A(Row1[113]), .Z(Output_2Row1[113]) );
  BUF_X4 U286 ( .A(Row1[190]), .Z(Output_2Row1[190]) );
  BUF_X4 U287 ( .A(Row1[189]), .Z(Output_2Row1[189]) );
  BUF_X4 U288 ( .A(Row1[125]), .Z(Output_2Row1[125]) );
  BUF_X4 U289 ( .A(Row1[191]), .Z(Output_2Row1[191]) );
  BUF_X4 U290 ( .A(Row1[64]), .Z(Output_2Row1[64]) );
  BUF_X4 U291 ( .A(Row1[65]), .Z(Output_2Row1[65]) );
  BUF_X4 U292 ( .A(Row1[66]), .Z(Output_2Row1[66]) );
  BUF_X4 U293 ( .A(Row1[67]), .Z(Output_2Row1[67]) );
  BUF_X4 U294 ( .A(Row1[68]), .Z(Output_2Row1[68]) );
  BUF_X4 U295 ( .A(Row1[69]), .Z(Output_2Row1[69]) );
  BUF_X4 U296 ( .A(Row1[70]), .Z(Output_2Row1[70]) );
  BUF_X4 U297 ( .A(Row1[71]), .Z(Output_2Row1[71]) );
  BUF_X4 U298 ( .A(Row1[72]), .Z(Output_2Row1[72]) );
  BUF_X4 U299 ( .A(Row1[73]), .Z(Output_2Row1[73]) );
  BUF_X4 U300 ( .A(Row1[74]), .Z(Output_2Row1[74]) );
  BUF_X4 U301 ( .A(Row1[80]), .Z(Output_2Row1[80]) );
  BUF_X4 U302 ( .A(Row1[81]), .Z(Output_2Row1[81]) );
  BUF_X4 U303 ( .A(Row1[82]), .Z(Output_2Row1[82]) );
  BUF_X4 U304 ( .A(Row1[83]), .Z(Output_2Row1[83]) );
  BUF_X4 U305 ( .A(Row1[84]), .Z(Output_2Row1[84]) );
  BUF_X4 U306 ( .A(Row1[85]), .Z(Output_2Row1[85]) );
  BUF_X4 U307 ( .A(Row1[86]), .Z(Output_2Row1[86]) );
  BUF_X4 U308 ( .A(Row1[87]), .Z(Output_2Row1[87]) );
  BUF_X4 U309 ( .A(Row1[88]), .Z(Output_2Row1[88]) );
  BUF_X4 U310 ( .A(Row1[89]), .Z(Output_2Row1[89]) );
  BUF_X4 U311 ( .A(Row1[90]), .Z(Output_2Row1[90]) );
  BUF_X4 U312 ( .A(Row1[96]), .Z(Output_2Row1[96]) );
  BUF_X4 U313 ( .A(Row1[97]), .Z(Output_2Row1[97]) );
  BUF_X4 U314 ( .A(Row1[98]), .Z(Output_2Row1[98]) );
  BUF_X4 U315 ( .A(Row1[99]), .Z(Output_2Row1[99]) );
  BUF_X4 U316 ( .A(Row1[100]), .Z(Output_2Row1[100]) );
  BUF_X4 U317 ( .A(Row1[101]), .Z(Output_2Row1[101]) );
  BUF_X4 U318 ( .A(Row1[102]), .Z(Output_2Row1[102]) );
  BUF_X4 U319 ( .A(Row1[103]), .Z(Output_2Row1[103]) );
  BUF_X4 U320 ( .A(Row1[104]), .Z(Output_2Row1[104]) );
  BUF_X4 U321 ( .A(Row1[105]), .Z(Output_2Row1[105]) );
  BUF_X4 U322 ( .A(Row1[106]), .Z(Output_2Row1[106]) );
  BUF_X4 U323 ( .A(Row1[246]), .Z(Output_2Row1[246]) );
  BUF_X4 U324 ( .A(Row1[247]), .Z(Output_2Row1[247]) );
  BUF_X4 U325 ( .A(Row1[243]), .Z(Output_2Row1[243]) );
  BUF_X4 U326 ( .A(Row1[240]), .Z(Output_2Row1[240]) );
  BUF_X4 U327 ( .A(Row1[245]), .Z(Output_2Row1[245]) );
  BUF_X4 U328 ( .A(Row1[244]), .Z(Output_2Row1[244]) );
  BUF_X4 U329 ( .A(Row1[242]), .Z(Output_2Row1[242]) );
  BUF_X4 U330 ( .A(Row1[241]), .Z(Output_2Row1[241]) );
  BUF_X4 U331 ( .A(Row1[254]), .Z(Output_2Row1[254]) );
  BUF_X4 U332 ( .A(Row1[253]), .Z(Output_2Row1[253]) );
  BUF_X4 U333 ( .A(Row1[255]), .Z(Output_2Row1[255]) );
  BUF_X4 U334 ( .A(Row1[254]), .Z(OutputCompute[254]) );
  BUF_X4 U335 ( .A(Row1[253]), .Z(OutputCompute[253]) );
  BUF_X4 U336 ( .A(Row1[255]), .Z(OutputCompute[255]) );
  BUF_X4 U337 ( .A(Row1[62]), .Z(OutputCompute[62]) );
  BUF_X4 U338 ( .A(Row1[61]), .Z(OutputCompute[61]) );
  BUF_X4 U339 ( .A(Row1[63]), .Z(OutputCompute[63]) );
  BUF_X4 U340 ( .A(Row1[126]), .Z(OutputCompute[126]) );
  BUF_X4 U341 ( .A(Row1[125]), .Z(OutputCompute[125]) );
  BUF_X4 U342 ( .A(Row1[127]), .Z(OutputCompute[127]) );
  BUF_X4 U343 ( .A(Row1[190]), .Z(OutputCompute[190]) );
  BUF_X4 U344 ( .A(Row1[189]), .Z(OutputCompute[189]) );
  BUF_X4 U345 ( .A(Row1[191]), .Z(OutputCompute[191]) );
  BUF_X4 U346 ( .A(PaddedRow[64]), .Z(WriteBus[64]) );
  BUF_X4 U347 ( .A(Row1[64]), .Z(OutputPaddedRow[64]) );
  BUF_X4 U348 ( .A(PaddedRow[65]), .Z(WriteBus[65]) );
  BUF_X4 U349 ( .A(Row1[65]), .Z(OutputPaddedRow[65]) );
  BUF_X4 U350 ( .A(PaddedRow[66]), .Z(WriteBus[66]) );
  BUF_X4 U351 ( .A(Row1[66]), .Z(OutputPaddedRow[66]) );
  BUF_X4 U352 ( .A(PaddedRow[67]), .Z(WriteBus[67]) );
  BUF_X4 U353 ( .A(Row1[67]), .Z(OutputPaddedRow[67]) );
  BUF_X4 U354 ( .A(PaddedRow[68]), .Z(WriteBus[68]) );
  BUF_X4 U355 ( .A(Row1[68]), .Z(OutputPaddedRow[68]) );
  BUF_X4 U356 ( .A(PaddedRow[69]), .Z(WriteBus[69]) );
  BUF_X4 U357 ( .A(Row1[69]), .Z(OutputPaddedRow[69]) );
  BUF_X4 U358 ( .A(PaddedRow[70]), .Z(WriteBus[70]) );
  BUF_X4 U359 ( .A(Row1[70]), .Z(OutputPaddedRow[70]) );
  BUF_X4 U360 ( .A(PaddedRow[71]), .Z(WriteBus[71]) );
  BUF_X4 U361 ( .A(Row1[71]), .Z(OutputPaddedRow[71]) );
  BUF_X4 U362 ( .A(PaddedRow[72]), .Z(WriteBus[72]) );
  BUF_X4 U363 ( .A(Row1[72]), .Z(OutputPaddedRow[72]) );
  BUF_X4 U364 ( .A(PaddedRow[73]), .Z(WriteBus[73]) );
  BUF_X4 U365 ( .A(Row1[73]), .Z(OutputPaddedRow[73]) );
  BUF_X4 U366 ( .A(PaddedRow[74]), .Z(WriteBus[74]) );
  BUF_X4 U367 ( .A(Row1[74]), .Z(OutputPaddedRow[74]) );
  BUF_X4 U368 ( .A(PaddedRow[80]), .Z(WriteBus[80]) );
  BUF_X4 U369 ( .A(Row1[80]), .Z(OutputPaddedRow[80]) );
  BUF_X4 U370 ( .A(PaddedRow[81]), .Z(WriteBus[81]) );
  BUF_X4 U371 ( .A(Row1[81]), .Z(OutputPaddedRow[81]) );
  BUF_X4 U372 ( .A(PaddedRow[82]), .Z(WriteBus[82]) );
  BUF_X4 U373 ( .A(Row1[82]), .Z(OutputPaddedRow[82]) );
  BUF_X4 U374 ( .A(PaddedRow[83]), .Z(WriteBus[83]) );
  BUF_X4 U375 ( .A(Row1[83]), .Z(OutputPaddedRow[83]) );
  BUF_X4 U376 ( .A(PaddedRow[84]), .Z(WriteBus[84]) );
  BUF_X4 U377 ( .A(Row1[84]), .Z(OutputPaddedRow[84]) );
  BUF_X4 U378 ( .A(PaddedRow[85]), .Z(WriteBus[85]) );
  BUF_X4 U379 ( .A(Row1[85]), .Z(OutputPaddedRow[85]) );
  BUF_X4 U380 ( .A(PaddedRow[86]), .Z(WriteBus[86]) );
  BUF_X4 U381 ( .A(Row1[86]), .Z(OutputPaddedRow[86]) );
  BUF_X4 U382 ( .A(PaddedRow[87]), .Z(WriteBus[87]) );
  BUF_X4 U383 ( .A(Row1[87]), .Z(OutputPaddedRow[87]) );
  BUF_X4 U384 ( .A(PaddedRow[88]), .Z(WriteBus[88]) );
  BUF_X4 U385 ( .A(Row1[88]), .Z(OutputPaddedRow[88]) );
  BUF_X4 U386 ( .A(PaddedRow[89]), .Z(WriteBus[89]) );
  BUF_X4 U387 ( .A(Row1[89]), .Z(OutputPaddedRow[89]) );
  BUF_X4 U388 ( .A(PaddedRow[100]), .Z(WriteBus[100]) );
  BUF_X4 U389 ( .A(Row1[100]), .Z(OutputPaddedRow[100]) );
  BUF_X4 U390 ( .A(PaddedRow[101]), .Z(WriteBus[101]) );
  BUF_X4 U391 ( .A(Row1[101]), .Z(OutputPaddedRow[101]) );
  BUF_X4 U392 ( .A(PaddedRow[102]), .Z(WriteBus[102]) );
  BUF_X4 U393 ( .A(Row1[102]), .Z(OutputPaddedRow[102]) );
  BUF_X4 U394 ( .A(PaddedRow[103]), .Z(WriteBus[103]) );
  BUF_X4 U395 ( .A(Row1[103]), .Z(OutputPaddedRow[103]) );
  BUF_X4 U396 ( .A(PaddedRow[104]), .Z(WriteBus[104]) );
  BUF_X4 U397 ( .A(Row1[104]), .Z(OutputPaddedRow[104]) );
  BUF_X4 U398 ( .A(PaddedRow[105]), .Z(WriteBus[105]) );
  BUF_X4 U399 ( .A(Row1[105]), .Z(OutputPaddedRow[105]) );
  BUF_X4 U400 ( .A(PaddedRow[106]), .Z(WriteBus[106]) );
  BUF_X4 U401 ( .A(Row1[106]), .Z(OutputPaddedRow[106]) );
  BUF_X4 U402 ( .A(PaddedRow[90]), .Z(WriteBus[90]) );
  BUF_X4 U403 ( .A(Row1[90]), .Z(OutputPaddedRow[90]) );
  BUF_X4 U404 ( .A(PaddedRow[96]), .Z(WriteBus[96]) );
  BUF_X4 U405 ( .A(Row1[96]), .Z(OutputPaddedRow[96]) );
  BUF_X4 U406 ( .A(PaddedRow[97]), .Z(WriteBus[97]) );
  BUF_X4 U407 ( .A(Row1[97]), .Z(OutputPaddedRow[97]) );
  BUF_X4 U408 ( .A(PaddedRow[98]), .Z(WriteBus[98]) );
  BUF_X4 U409 ( .A(Row1[98]), .Z(OutputPaddedRow[98]) );
  BUF_X4 U410 ( .A(PaddedRow[99]), .Z(WriteBus[99]) );
  BUF_X4 U411 ( .A(Row1[99]), .Z(OutputPaddedRow[99]) );
  INV_X4 U412 ( .A(n2960), .ZN(n4800) );
  BUF_X4 U413 ( .A(Row1[60]), .Z(OutputCompute[60]) );
  BUF_X4 U414 ( .A(Row1[188]), .Z(OutputCompute[188]) );
  BUF_X4 U415 ( .A(Row1[124]), .Z(OutputCompute[124]) );
  BUF_X4 U416 ( .A(Row1[252]), .Z(OutputCompute[252]) );
  BUF_X4 U417 ( .A(Row1[96]), .Z(Output_1Row1[96]) );
  BUF_X4 U418 ( .A(Row1[112]), .Z(Output_1Row1[112]) );
  BUF_X4 U419 ( .A(Row1[64]), .Z(Output_1Row1[64]) );
  BUF_X4 U420 ( .A(Row1[80]), .Z(Output_1Row1[80]) );
  BUF_X4 U421 ( .A(Row1[73]), .Z(Output_1Row1[73]) );
  BUF_X4 U422 ( .A(Row1[89]), .Z(Output_1Row1[89]) );
  BUF_X4 U423 ( .A(Row1[72]), .Z(Output_1Row1[72]) );
  BUF_X4 U424 ( .A(Row1[88]), .Z(Output_1Row1[88]) );
  BUF_X4 U425 ( .A(Row1[71]), .Z(Output_1Row1[71]) );
  BUF_X4 U426 ( .A(Row1[87]), .Z(Output_1Row1[87]) );
  BUF_X4 U427 ( .A(Row1[70]), .Z(Output_1Row1[70]) );
  BUF_X4 U428 ( .A(Row1[86]), .Z(Output_1Row1[86]) );
  BUF_X4 U429 ( .A(Row1[69]), .Z(Output_1Row1[69]) );
  BUF_X4 U430 ( .A(Row1[85]), .Z(Output_1Row1[85]) );
  BUF_X4 U431 ( .A(Row1[68]), .Z(Output_1Row1[68]) );
  BUF_X4 U432 ( .A(Row1[84]), .Z(Output_1Row1[84]) );
  BUF_X4 U433 ( .A(Row1[67]), .Z(Output_1Row1[67]) );
  BUF_X4 U434 ( .A(Row1[83]), .Z(Output_1Row1[83]) );
  BUF_X4 U435 ( .A(Row1[66]), .Z(Output_1Row1[66]) );
  BUF_X4 U436 ( .A(Row1[82]), .Z(Output_1Row1[82]) );
  BUF_X4 U437 ( .A(Row1[65]), .Z(Output_1Row1[65]) );
  BUF_X4 U438 ( .A(Row1[81]), .Z(Output_1Row1[81]) );
  BUF_X4 U439 ( .A(Row1[105]), .Z(Output_1Row1[105]) );
  BUF_X4 U440 ( .A(Row1[121]), .Z(Output_1Row1[121]) );
  BUF_X4 U441 ( .A(Row1[104]), .Z(Output_1Row1[104]) );
  BUF_X4 U442 ( .A(Row1[120]), .Z(Output_1Row1[120]) );
  BUF_X4 U443 ( .A(Row1[103]), .Z(Output_1Row1[103]) );
  BUF_X4 U444 ( .A(Row1[119]), .Z(Output_1Row1[119]) );
  BUF_X4 U445 ( .A(Row1[102]), .Z(Output_1Row1[102]) );
  BUF_X4 U446 ( .A(Row1[118]), .Z(Output_1Row1[118]) );
  BUF_X4 U447 ( .A(Row1[101]), .Z(Output_1Row1[101]) );
  BUF_X4 U448 ( .A(Row1[117]), .Z(Output_1Row1[117]) );
  BUF_X4 U449 ( .A(Row1[100]), .Z(Output_1Row1[100]) );
  BUF_X4 U450 ( .A(Row1[116]), .Z(Output_1Row1[116]) );
  BUF_X4 U451 ( .A(Row1[99]), .Z(Output_1Row1[99]) );
  BUF_X4 U452 ( .A(Row1[115]), .Z(Output_1Row1[115]) );
  BUF_X4 U453 ( .A(Row1[98]), .Z(Output_1Row1[98]) );
  BUF_X4 U454 ( .A(Row1[114]), .Z(Output_1Row1[114]) );
  BUF_X4 U455 ( .A(Row1[97]), .Z(Output_1Row1[97]) );
  BUF_X4 U456 ( .A(Row1[113]), .Z(Output_1Row1[113]) );
  BUF_X4 U457 ( .A(PaddedRow[48]), .Z(WriteBus[48]) );
  BUF_X4 U458 ( .A(Row1[48]), .Z(OutputPaddedRow[48]) );
  BUF_X4 U459 ( .A(PaddedRow[49]), .Z(WriteBus[49]) );
  BUF_X4 U460 ( .A(Row1[49]), .Z(OutputPaddedRow[49]) );
  BUF_X4 U461 ( .A(PaddedRow[50]), .Z(WriteBus[50]) );
  BUF_X4 U462 ( .A(Row1[50]), .Z(OutputPaddedRow[50]) );
  BUF_X4 U463 ( .A(PaddedRow[51]), .Z(WriteBus[51]) );
  BUF_X4 U464 ( .A(Row1[51]), .Z(OutputPaddedRow[51]) );
  BUF_X4 U465 ( .A(PaddedRow[52]), .Z(WriteBus[52]) );
  BUF_X4 U466 ( .A(Row1[52]), .Z(OutputPaddedRow[52]) );
  BUF_X4 U467 ( .A(PaddedRow[53]), .Z(WriteBus[53]) );
  BUF_X4 U468 ( .A(Row1[53]), .Z(OutputPaddedRow[53]) );
  BUF_X4 U469 ( .A(PaddedRow[54]), .Z(WriteBus[54]) );
  BUF_X4 U470 ( .A(Row1[54]), .Z(OutputPaddedRow[54]) );
  BUF_X4 U471 ( .A(PaddedRow[55]), .Z(WriteBus[55]) );
  BUF_X4 U472 ( .A(Row1[55]), .Z(OutputPaddedRow[55]) );
  BUF_X4 U473 ( .A(PaddedRow[56]), .Z(WriteBus[56]) );
  BUF_X4 U474 ( .A(Row1[56]), .Z(OutputPaddedRow[56]) );
  BUF_X4 U475 ( .A(PaddedRow[57]), .Z(WriteBus[57]) );
  BUF_X4 U476 ( .A(Row1[57]), .Z(OutputPaddedRow[57]) );
  BUF_X4 U477 ( .A(PaddedRow[58]), .Z(WriteBus[58]) );
  BUF_X4 U478 ( .A(Row1[58]), .Z(OutputPaddedRow[58]) );
  BUF_X4 U479 ( .A(PaddedRow[59]), .Z(WriteBus[59]) );
  BUF_X4 U480 ( .A(Row1[59]), .Z(OutputPaddedRow[59]) );
  BUF_X4 U481 ( .A(PaddedRow[60]), .Z(WriteBus[60]) );
  BUF_X4 U482 ( .A(Row1[60]), .Z(OutputPaddedRow[60]) );
  BUF_X4 U483 ( .A(PaddedRow[61]), .Z(WriteBus[61]) );
  BUF_X4 U484 ( .A(Row1[61]), .Z(OutputPaddedRow[61]) );
  BUF_X4 U485 ( .A(PaddedRow[62]), .Z(WriteBus[62]) );
  BUF_X4 U486 ( .A(Row1[62]), .Z(OutputPaddedRow[62]) );
  BUF_X4 U487 ( .A(PaddedRow[63]), .Z(WriteBus[63]) );
  BUF_X4 U488 ( .A(Row1[63]), .Z(OutputPaddedRow[63]) );
  BUF_X4 U489 ( .A(PaddedRow[112]), .Z(WriteBus[112]) );
  BUF_X4 U490 ( .A(Row1[112]), .Z(OutputPaddedRow[112]) );
  BUF_X4 U491 ( .A(PaddedRow[113]), .Z(WriteBus[113]) );
  BUF_X4 U492 ( .A(Row1[113]), .Z(OutputPaddedRow[113]) );
  BUF_X4 U493 ( .A(PaddedRow[114]), .Z(WriteBus[114]) );
  BUF_X4 U494 ( .A(Row1[114]), .Z(OutputPaddedRow[114]) );
  BUF_X4 U495 ( .A(PaddedRow[115]), .Z(WriteBus[115]) );
  BUF_X4 U496 ( .A(Row1[115]), .Z(OutputPaddedRow[115]) );
  BUF_X4 U497 ( .A(PaddedRow[116]), .Z(WriteBus[116]) );
  BUF_X4 U498 ( .A(Row1[116]), .Z(OutputPaddedRow[116]) );
  BUF_X4 U499 ( .A(PaddedRow[117]), .Z(WriteBus[117]) );
  BUF_X4 U500 ( .A(Row1[117]), .Z(OutputPaddedRow[117]) );
  BUF_X4 U501 ( .A(PaddedRow[118]), .Z(WriteBus[118]) );
  BUF_X4 U502 ( .A(Row1[118]), .Z(OutputPaddedRow[118]) );
  BUF_X4 U503 ( .A(PaddedRow[119]), .Z(WriteBus[119]) );
  BUF_X4 U504 ( .A(Row1[119]), .Z(OutputPaddedRow[119]) );
  BUF_X4 U505 ( .A(PaddedRow[120]), .Z(WriteBus[120]) );
  BUF_X4 U506 ( .A(Row1[120]), .Z(OutputPaddedRow[120]) );
  BUF_X4 U507 ( .A(PaddedRow[121]), .Z(WriteBus[121]) );
  BUF_X4 U508 ( .A(Row1[121]), .Z(OutputPaddedRow[121]) );
  BUF_X4 U509 ( .A(PaddedRow[122]), .Z(WriteBus[122]) );
  BUF_X4 U510 ( .A(Row1[122]), .Z(OutputPaddedRow[122]) );
  BUF_X4 U511 ( .A(PaddedRow[123]), .Z(WriteBus[123]) );
  BUF_X4 U512 ( .A(Row1[123]), .Z(OutputPaddedRow[123]) );
  BUF_X4 U513 ( .A(PaddedRow[124]), .Z(WriteBus[124]) );
  BUF_X4 U514 ( .A(Row1[124]), .Z(OutputPaddedRow[124]) );
  BUF_X4 U515 ( .A(PaddedRow[125]), .Z(WriteBus[125]) );
  BUF_X4 U516 ( .A(Row1[125]), .Z(OutputPaddedRow[125]) );
  BUF_X4 U517 ( .A(PaddedRow[126]), .Z(WriteBus[126]) );
  BUF_X4 U518 ( .A(Row1[126]), .Z(OutputPaddedRow[126]) );
  BUF_X4 U519 ( .A(PaddedRow[127]), .Z(WriteBus[127]) );
  BUF_X4 U520 ( .A(Row1[127]), .Z(OutputPaddedRow[127]) );
  BUF_X4 U521 ( .A(PaddedRow[176]), .Z(WriteBus[176]) );
  BUF_X4 U522 ( .A(Row1[176]), .Z(OutputPaddedRow[176]) );
  BUF_X4 U523 ( .A(PaddedRow[177]), .Z(WriteBus[177]) );
  BUF_X4 U524 ( .A(Row1[177]), .Z(OutputPaddedRow[177]) );
  BUF_X4 U525 ( .A(PaddedRow[178]), .Z(WriteBus[178]) );
  BUF_X4 U526 ( .A(Row1[178]), .Z(OutputPaddedRow[178]) );
  BUF_X4 U527 ( .A(PaddedRow[179]), .Z(WriteBus[179]) );
  BUF_X4 U528 ( .A(Row1[179]), .Z(OutputPaddedRow[179]) );
  BUF_X4 U529 ( .A(PaddedRow[180]), .Z(WriteBus[180]) );
  BUF_X4 U530 ( .A(Row1[180]), .Z(OutputPaddedRow[180]) );
  BUF_X4 U531 ( .A(PaddedRow[181]), .Z(WriteBus[181]) );
  BUF_X4 U532 ( .A(Row1[181]), .Z(OutputPaddedRow[181]) );
  BUF_X4 U533 ( .A(PaddedRow[182]), .Z(WriteBus[182]) );
  BUF_X4 U534 ( .A(Row1[182]), .Z(OutputPaddedRow[182]) );
  BUF_X4 U535 ( .A(PaddedRow[183]), .Z(WriteBus[183]) );
  BUF_X4 U536 ( .A(Row1[183]), .Z(OutputPaddedRow[183]) );
  BUF_X4 U537 ( .A(PaddedRow[184]), .Z(WriteBus[184]) );
  BUF_X4 U538 ( .A(Row1[184]), .Z(OutputPaddedRow[184]) );
  BUF_X4 U539 ( .A(PaddedRow[185]), .Z(WriteBus[185]) );
  BUF_X4 U540 ( .A(Row1[185]), .Z(OutputPaddedRow[185]) );
  BUF_X4 U541 ( .A(PaddedRow[186]), .Z(WriteBus[186]) );
  BUF_X4 U542 ( .A(Row1[186]), .Z(OutputPaddedRow[186]) );
  BUF_X4 U543 ( .A(PaddedRow[187]), .Z(WriteBus[187]) );
  BUF_X4 U544 ( .A(Row1[187]), .Z(OutputPaddedRow[187]) );
  BUF_X4 U545 ( .A(PaddedRow[188]), .Z(WriteBus[188]) );
  BUF_X4 U546 ( .A(Row1[188]), .Z(OutputPaddedRow[188]) );
  BUF_X4 U547 ( .A(PaddedRow[189]), .Z(WriteBus[189]) );
  BUF_X4 U548 ( .A(Row1[189]), .Z(OutputPaddedRow[189]) );
  BUF_X4 U549 ( .A(PaddedRow[190]), .Z(WriteBus[190]) );
  BUF_X4 U550 ( .A(Row1[190]), .Z(OutputPaddedRow[190]) );
  BUF_X4 U551 ( .A(PaddedRow[191]), .Z(WriteBus[191]) );
  BUF_X4 U552 ( .A(Row1[191]), .Z(OutputPaddedRow[191]) );
  BUF_X4 U553 ( .A(PaddedRow[240]), .Z(WriteBus[240]) );
  BUF_X4 U554 ( .A(Row1[240]), .Z(OutputPaddedRow[240]) );
  BUF_X4 U555 ( .A(PaddedRow[241]), .Z(WriteBus[241]) );
  BUF_X4 U556 ( .A(Row1[241]), .Z(OutputPaddedRow[241]) );
  BUF_X4 U557 ( .A(PaddedRow[242]), .Z(WriteBus[242]) );
  BUF_X4 U558 ( .A(Row1[242]), .Z(OutputPaddedRow[242]) );
  BUF_X4 U559 ( .A(PaddedRow[243]), .Z(WriteBus[243]) );
  BUF_X4 U560 ( .A(Row1[243]), .Z(OutputPaddedRow[243]) );
  BUF_X4 U561 ( .A(PaddedRow[244]), .Z(WriteBus[244]) );
  BUF_X4 U562 ( .A(Row1[244]), .Z(OutputPaddedRow[244]) );
  BUF_X4 U563 ( .A(PaddedRow[245]), .Z(WriteBus[245]) );
  BUF_X4 U564 ( .A(Row1[245]), .Z(OutputPaddedRow[245]) );
  BUF_X4 U565 ( .A(PaddedRow[246]), .Z(WriteBus[246]) );
  BUF_X4 U566 ( .A(Row1[246]), .Z(OutputPaddedRow[246]) );
  BUF_X4 U567 ( .A(PaddedRow[247]), .Z(WriteBus[247]) );
  BUF_X4 U568 ( .A(Row1[247]), .Z(OutputPaddedRow[247]) );
  BUF_X4 U569 ( .A(PaddedRow[248]), .Z(WriteBus[248]) );
  BUF_X4 U570 ( .A(Row1[248]), .Z(OutputPaddedRow[248]) );
  BUF_X4 U571 ( .A(PaddedRow[249]), .Z(WriteBus[249]) );
  BUF_X4 U572 ( .A(Row1[249]), .Z(OutputPaddedRow[249]) );
  BUF_X4 U573 ( .A(PaddedRow[250]), .Z(WriteBus[250]) );
  BUF_X4 U574 ( .A(Row1[250]), .Z(OutputPaddedRow[250]) );
  BUF_X4 U575 ( .A(PaddedRow[251]), .Z(WriteBus[251]) );
  BUF_X4 U576 ( .A(Row1[251]), .Z(OutputPaddedRow[251]) );
  BUF_X4 U577 ( .A(PaddedRow[252]), .Z(WriteBus[252]) );
  BUF_X4 U578 ( .A(Row1[252]), .Z(OutputPaddedRow[252]) );
  BUF_X4 U579 ( .A(PaddedRow[253]), .Z(WriteBus[253]) );
  BUF_X4 U580 ( .A(Row1[253]), .Z(OutputPaddedRow[253]) );
  BUF_X4 U581 ( .A(PaddedRow[254]), .Z(WriteBus[254]) );
  BUF_X4 U582 ( .A(Row1[254]), .Z(OutputPaddedRow[254]) );
  BUF_X4 U583 ( .A(PaddedRow[255]), .Z(WriteBus[255]) );
  BUF_X4 U584 ( .A(Row1[255]), .Z(OutputPaddedRow[255]) );
  BUF_X4 U585 ( .A(Row1[248]), .Z(OutputCompute[248]) );
  BUF_X4 U586 ( .A(Row1[250]), .Z(OutputCompute[250]) );
  BUF_X4 U587 ( .A(Row1[184]), .Z(OutputCompute[184]) );
  BUF_X4 U588 ( .A(Row1[249]), .Z(OutputCompute[249]) );
  BUF_X4 U589 ( .A(Row1[186]), .Z(OutputCompute[186]) );
  BUF_X4 U590 ( .A(Row1[185]), .Z(OutputCompute[185]) );
  BUF_X4 U591 ( .A(Row1[120]), .Z(OutputCompute[120]) );
  BUF_X4 U592 ( .A(Row1[122]), .Z(OutputCompute[122]) );
  BUF_X4 U593 ( .A(Row1[121]), .Z(OutputCompute[121]) );
  BUF_X4 U594 ( .A(Row1[56]), .Z(OutputCompute[56]) );
  BUF_X4 U595 ( .A(Row1[58]), .Z(OutputCompute[58]) );
  BUF_X4 U596 ( .A(Row1[57]), .Z(OutputCompute[57]) );
  BUF_X4 U597 ( .A(Row1[251]), .Z(OutputCompute[251]) );
  BUF_X4 U598 ( .A(Row1[123]), .Z(OutputCompute[123]) );
  BUF_X4 U599 ( .A(Row1[187]), .Z(OutputCompute[187]) );
  BUF_X4 U600 ( .A(Row1[59]), .Z(OutputCompute[59]) );
  BUF_X4 U601 ( .A(Row1[249]), .Z(Output_1Row1[249]) );
  BUF_X4 U602 ( .A(Row1[248]), .Z(Output_1Row1[248]) );
  BUF_X4 U603 ( .A(Row1[247]), .Z(Output_1Row1[247]) );
  BUF_X4 U604 ( .A(Row1[246]), .Z(Output_1Row1[246]) );
  BUF_X4 U605 ( .A(Row1[245]), .Z(Output_1Row1[245]) );
  BUF_X4 U606 ( .A(Row1[244]), .Z(Output_1Row1[244]) );
  BUF_X4 U607 ( .A(Row1[243]), .Z(Output_1Row1[243]) );
  BUF_X4 U608 ( .A(Row1[242]), .Z(Output_1Row1[242]) );
  BUF_X4 U609 ( .A(Row1[241]), .Z(Output_1Row1[241]) );
  OAI21_X2 U610 ( .B1(reset), .B2(n37), .A(n38), .ZN(\U4/Z_3 ) );
  NOR2_X2 U611 ( .A1(n51), .A2(n4768), .ZN(n85) );
  AOI21_X2 U612 ( .B1(n4768), .B2(n42), .A(n1830), .ZN(\U3/U1/Z_0 ) );
  NOR2_X2 U613 ( .A1(n56), .A2(n4770), .ZN(n81) );
  INV_X4 U614 ( .A(n56), .ZN(n4798) );
  INV_X4 U615 ( .A(n55), .ZN(n4802) );
  INV_X4 U616 ( .A(n42), .ZN(n4801) );
  BUF_X4 U617 ( .A(Row1[64]), .Z(OutputCompute[64]) );
  BUF_X4 U618 ( .A(Row1[65]), .Z(OutputCompute[65]) );
  BUF_X4 U619 ( .A(Row1[66]), .Z(OutputCompute[66]) );
  BUF_X4 U620 ( .A(Row1[67]), .Z(OutputCompute[67]) );
  BUF_X4 U621 ( .A(Row1[68]), .Z(OutputCompute[68]) );
  BUF_X4 U622 ( .A(Row1[69]), .Z(OutputCompute[69]) );
  BUF_X4 U623 ( .A(Row1[70]), .Z(OutputCompute[70]) );
  BUF_X4 U624 ( .A(Row1[71]), .Z(OutputCompute[71]) );
  BUF_X4 U625 ( .A(Row1[72]), .Z(OutputCompute[72]) );
  BUF_X4 U626 ( .A(Row1[73]), .Z(OutputCompute[73]) );
  BUF_X4 U627 ( .A(Row1[74]), .Z(OutputCompute[74]) );
  BUF_X4 U628 ( .A(Row1[80]), .Z(OutputCompute[80]) );
  BUF_X4 U629 ( .A(Row1[81]), .Z(OutputCompute[81]) );
  BUF_X4 U630 ( .A(Row1[82]), .Z(OutputCompute[82]) );
  BUF_X4 U631 ( .A(Row1[83]), .Z(OutputCompute[83]) );
  BUF_X4 U632 ( .A(Row1[84]), .Z(OutputCompute[84]) );
  BUF_X4 U633 ( .A(Row1[85]), .Z(OutputCompute[85]) );
  BUF_X4 U634 ( .A(Row1[86]), .Z(OutputCompute[86]) );
  BUF_X4 U635 ( .A(Row1[87]), .Z(OutputCompute[87]) );
  BUF_X4 U636 ( .A(Row1[88]), .Z(OutputCompute[88]) );
  BUF_X4 U637 ( .A(Row1[89]), .Z(OutputCompute[89]) );
  BUF_X4 U638 ( .A(Row1[90]), .Z(OutputCompute[90]) );
  BUF_X4 U639 ( .A(Row1[96]), .Z(OutputCompute[96]) );
  BUF_X4 U640 ( .A(Row1[97]), .Z(OutputCompute[97]) );
  BUF_X4 U641 ( .A(Row1[98]), .Z(OutputCompute[98]) );
  BUF_X4 U642 ( .A(Row1[99]), .Z(OutputCompute[99]) );
  BUF_X4 U643 ( .A(Row1[100]), .Z(OutputCompute[100]) );
  BUF_X4 U644 ( .A(Row1[101]), .Z(OutputCompute[101]) );
  BUF_X4 U645 ( .A(Row1[102]), .Z(OutputCompute[102]) );
  BUF_X4 U646 ( .A(Row1[103]), .Z(OutputCompute[103]) );
  BUF_X4 U647 ( .A(Row1[104]), .Z(OutputCompute[104]) );
  BUF_X4 U648 ( .A(Row1[105]), .Z(OutputCompute[105]) );
  BUF_X4 U649 ( .A(Row1[106]), .Z(OutputCompute[106]) );
  BUF_X4 U650 ( .A(Row1[112]), .Z(OutputCompute[112]) );
  BUF_X4 U651 ( .A(Row1[113]), .Z(OutputCompute[113]) );
  BUF_X4 U652 ( .A(Row1[114]), .Z(OutputCompute[114]) );
  BUF_X4 U653 ( .A(Row1[115]), .Z(OutputCompute[115]) );
  BUF_X4 U654 ( .A(Row1[116]), .Z(OutputCompute[116]) );
  BUF_X4 U655 ( .A(Row1[117]), .Z(OutputCompute[117]) );
  BUF_X4 U656 ( .A(Row1[118]), .Z(OutputCompute[118]) );
  BUF_X4 U657 ( .A(Row1[119]), .Z(OutputCompute[119]) );
  BUF_X4 U658 ( .A(Row1[48]), .Z(OutputCompute[48]) );
  BUF_X4 U659 ( .A(Row1[49]), .Z(OutputCompute[49]) );
  BUF_X4 U660 ( .A(Row1[50]), .Z(OutputCompute[50]) );
  BUF_X4 U661 ( .A(Row1[51]), .Z(OutputCompute[51]) );
  BUF_X4 U662 ( .A(Row1[52]), .Z(OutputCompute[52]) );
  BUF_X4 U663 ( .A(Row1[53]), .Z(OutputCompute[53]) );
  BUF_X4 U664 ( .A(Row1[54]), .Z(OutputCompute[54]) );
  BUF_X4 U665 ( .A(Row1[55]), .Z(OutputCompute[55]) );
  BUF_X4 U666 ( .A(Row1[240]), .Z(OutputCompute[240]) );
  BUF_X4 U667 ( .A(Row1[241]), .Z(OutputCompute[241]) );
  BUF_X4 U668 ( .A(Row1[242]), .Z(OutputCompute[242]) );
  BUF_X4 U669 ( .A(Row1[243]), .Z(OutputCompute[243]) );
  BUF_X4 U670 ( .A(Row1[244]), .Z(OutputCompute[244]) );
  BUF_X4 U671 ( .A(Row1[245]), .Z(OutputCompute[245]) );
  BUF_X4 U672 ( .A(Row1[246]), .Z(OutputCompute[246]) );
  BUF_X4 U673 ( .A(Row1[247]), .Z(OutputCompute[247]) );
  BUF_X4 U674 ( .A(Row1[74]), .Z(Output_1Row1[74]) );
  BUF_X4 U675 ( .A(Row1[106]), .Z(Output_1Row1[106]) );
  BUF_X4 U676 ( .A(Row1[250]), .Z(Output_1Row1[250]) );
  BUF_X4 U677 ( .A(Row1[90]), .Z(Output_1Row1[90]) );
  BUF_X4 U678 ( .A(Row1[122]), .Z(Output_1Row1[122]) );
  BUF_X4 U679 ( .A(\U3/U9/Z_0 ), .Z(ArbiterPos[2]) );
  BUF_X4 U680 ( .A(\U3/U9/Z_1 ), .Z(ArbiterPos[3]) );
  BUF_X4 U681 ( .A(\U3/U9/Z_2 ), .Z(ArbiterPos[4]) );
  BUF_X4 U682 ( .A(\U3/U9/Z_3 ), .Z(ArbiterPos[5]) );
  BUF_X4 U683 ( .A(\U3/U9/Z_4 ), .Z(ArbiterPos[6]) );
  BUF_X4 U684 ( .A(\U3/U9/Z_5 ), .Z(ArbiterPos[7]) );
  BUF_X4 U685 ( .A(\U3/U9/Z_6 ), .Z(ArbiterPos[8]) );
  BUF_X4 U686 ( .A(\U3/U9/Z_7 ), .Z(ArbiterPos[9]) );
  BUF_X4 U687 ( .A(\U3/U9/Z_8 ), .Z(ArbiterPos[10]) );
  BUF_X4 U688 ( .A(\U3/U9/Z_9 ), .Z(ArbiterPos[11]) );
  BUF_X4 U689 ( .A(\U3/U9/Z_10 ), .Z(ArbiterPos[12]) );
  BUF_X4 U690 ( .A(Row1[59]), .Z(Output_1Row1[59]) );
  BUF_X4 U691 ( .A(Row1[60]), .Z(Output_1Row1[60]) );
  BUF_X4 U692 ( .A(Row1[61]), .Z(Output_1Row1[61]) );
  BUF_X4 U693 ( .A(Row1[62]), .Z(Output_1Row1[62]) );
  BUF_X4 U694 ( .A(Row1[63]), .Z(Output_1Row1[63]) );
  BUF_X4 U695 ( .A(Row1[123]), .Z(Output_1Row1[123]) );
  BUF_X4 U696 ( .A(Row1[124]), .Z(Output_1Row1[124]) );
  BUF_X4 U697 ( .A(Row1[125]), .Z(Output_1Row1[125]) );
  BUF_X4 U698 ( .A(Row1[126]), .Z(Output_1Row1[126]) );
  BUF_X4 U699 ( .A(Row1[127]), .Z(Output_1Row1[127]) );
  BUF_X4 U700 ( .A(Row1[187]), .Z(Output_1Row1[187]) );
  BUF_X4 U701 ( .A(Row1[188]), .Z(Output_1Row1[188]) );
  BUF_X4 U702 ( .A(Row1[189]), .Z(Output_1Row1[189]) );
  BUF_X4 U703 ( .A(Row1[190]), .Z(Output_1Row1[190]) );
  BUF_X4 U704 ( .A(Row1[191]), .Z(Output_1Row1[191]) );
  BUF_X4 U705 ( .A(Row1[251]), .Z(Output_1Row1[251]) );
  BUF_X4 U706 ( .A(Row1[252]), .Z(Output_1Row1[252]) );
  BUF_X4 U707 ( .A(Row1[253]), .Z(Output_1Row1[253]) );
  BUF_X4 U708 ( .A(Row1[254]), .Z(Output_1Row1[254]) );
  BUF_X4 U709 ( .A(Row1[255]), .Z(Output_1Row1[255]) );
  BUF_X4 U710 ( .A(Row1[57]), .Z(Output_2Row1[57]) );
  BUF_X4 U711 ( .A(Row1[59]), .Z(Output_2Row1[59]) );
  BUF_X4 U712 ( .A(Row1[123]), .Z(Output_2Row1[123]) );
  BUF_X4 U713 ( .A(Row1[58]), .Z(Output_2Row1[58]) );
  BUF_X4 U714 ( .A(Row1[122]), .Z(Output_2Row1[122]) );
  BUF_X4 U715 ( .A(Row1[56]), .Z(Output_2Row1[56]) );
  BUF_X4 U716 ( .A(Row1[60]), .Z(Output_2Row1[60]) );
  BUF_X4 U717 ( .A(Row1[120]), .Z(Output_2Row1[120]) );
  BUF_X4 U718 ( .A(Row1[124]), .Z(Output_2Row1[124]) );
  BUF_X4 U719 ( .A(Row1[184]), .Z(Output_2Row1[184]) );
  BUF_X4 U720 ( .A(Row1[188]), .Z(Output_2Row1[188]) );
  BUF_X4 U721 ( .A(Row1[121]), .Z(Output_2Row1[121]) );
  BUF_X4 U722 ( .A(Row1[185]), .Z(Output_2Row1[185]) );
  BUF_X4 U723 ( .A(Row1[186]), .Z(Output_2Row1[186]) );
  BUF_X4 U724 ( .A(Row1[187]), .Z(Output_2Row1[187]) );
  BUF_X4 U725 ( .A(Row2[56]), .Z(Output_2Row2[56]) );
  BUF_X4 U726 ( .A(Row2[60]), .Z(Output_2Row2[60]) );
  BUF_X4 U727 ( .A(Row2[120]), .Z(Output_2Row2[120]) );
  BUF_X4 U728 ( .A(Row2[124]), .Z(Output_2Row2[124]) );
  BUF_X4 U729 ( .A(Row2[184]), .Z(Output_2Row2[184]) );
  BUF_X4 U730 ( .A(Row2[188]), .Z(Output_2Row2[188]) );
  BUF_X4 U731 ( .A(Row1[248]), .Z(Output_2Row1[248]) );
  BUF_X4 U732 ( .A(Row1[252]), .Z(Output_2Row1[252]) );
  BUF_X4 U733 ( .A(Row2[185]), .Z(Output_2Row2[185]) );
  BUF_X4 U734 ( .A(Row1[249]), .Z(Output_2Row1[249]) );
  BUF_X4 U735 ( .A(Row2[58]), .Z(Output_2Row2[58]) );
  BUF_X4 U736 ( .A(Row2[122]), .Z(Output_2Row2[122]) );
  BUF_X4 U737 ( .A(Row2[186]), .Z(Output_2Row2[186]) );
  BUF_X4 U738 ( .A(Row1[250]), .Z(Output_2Row1[250]) );
  BUF_X4 U739 ( .A(Row2[59]), .Z(Output_2Row2[59]) );
  BUF_X4 U740 ( .A(Row2[123]), .Z(Output_2Row2[123]) );
  BUF_X4 U741 ( .A(Row2[187]), .Z(Output_2Row2[187]) );
  BUF_X4 U742 ( .A(Row1[251]), .Z(Output_2Row1[251]) );
  BUF_X4 U743 ( .A(Row2[54]), .Z(Output_2Row2[54]) );
  BUF_X4 U744 ( .A(Row2[55]), .Z(Output_2Row2[55]) );
  BUF_X4 U745 ( .A(Row2[182]), .Z(Output_2Row2[182]) );
  BUF_X4 U746 ( .A(Row2[183]), .Z(Output_2Row2[183]) );
  BUF_X4 U747 ( .A(Row2[118]), .Z(Output_2Row2[118]) );
  BUF_X4 U748 ( .A(Row2[119]), .Z(Output_2Row2[119]) );
  BUF_X4 U749 ( .A(Row2[48]), .Z(Output_2Row2[48]) );
  BUF_X4 U750 ( .A(Row2[50]), .Z(Output_2Row2[50]) );
  BUF_X4 U751 ( .A(Row2[49]), .Z(Output_2Row2[49]) );
  BUF_X4 U752 ( .A(Row2[51]), .Z(Output_2Row2[51]) );
  BUF_X4 U753 ( .A(Row2[53]), .Z(Output_2Row2[53]) );
  BUF_X4 U754 ( .A(Row2[52]), .Z(Output_2Row2[52]) );
  BUF_X4 U755 ( .A(Row2[179]), .Z(Output_2Row2[179]) );
  BUF_X4 U756 ( .A(Row2[181]), .Z(Output_2Row2[181]) );
  BUF_X4 U757 ( .A(Row2[180]), .Z(Output_2Row2[180]) );
  BUF_X4 U758 ( .A(Row2[115]), .Z(Output_2Row2[115]) );
  BUF_X4 U759 ( .A(Row2[112]), .Z(Output_2Row2[112]) );
  BUF_X4 U760 ( .A(Row2[117]), .Z(Output_2Row2[117]) );
  BUF_X4 U761 ( .A(Row2[116]), .Z(Output_2Row2[116]) );
  BUF_X4 U762 ( .A(Row2[178]), .Z(Output_2Row2[178]) );
  BUF_X4 U763 ( .A(Row2[177]), .Z(Output_2Row2[177]) );
  BUF_X4 U764 ( .A(Row2[176]), .Z(Output_2Row2[176]) );
  BUF_X4 U765 ( .A(Row2[114]), .Z(Output_2Row2[114]) );
  BUF_X4 U766 ( .A(Row2[113]), .Z(Output_2Row2[113]) );
  BUF_X4 U767 ( .A(Row2[62]), .Z(Output_2Row2[62]) );
  BUF_X4 U768 ( .A(Row2[190]), .Z(Output_2Row2[190]) );
  BUF_X4 U769 ( .A(Row2[126]), .Z(Output_2Row2[126]) );
  BUF_X4 U770 ( .A(Row2[61]), .Z(Output_2Row2[61]) );
  BUF_X4 U771 ( .A(Row2[189]), .Z(Output_2Row2[189]) );
  BUF_X4 U772 ( .A(Row2[125]), .Z(Output_2Row2[125]) );
  BUF_X4 U773 ( .A(Row2[63]), .Z(Output_2Row2[63]) );
  BUF_X4 U774 ( .A(Row2[191]), .Z(Output_2Row2[191]) );
  BUF_X4 U775 ( .A(Row2[127]), .Z(Output_2Row2[127]) );
  BUF_X4 U776 ( .A(Row2[57]), .Z(Output_2Row2[57]) );
  BUF_X4 U777 ( .A(Row2[121]), .Z(Output_2Row2[121]) );
  AOI22_X2 U778 ( .A1(\U3/U8/DATA2_1 ), .A2(n4799), .B1(\U3/U8/DATA1_1 ), .B2(
        n4768), .ZN(n76) );
  AOI22_X2 U779 ( .A1(\U3/U8/DATA2_0 ), .A2(n4799), .B1(\U3/U8/DATA1_0 ), .B2(
        n4768), .ZN(n77) );
  BUF_X4 U780 ( .A(Row1[176]), .Z(OutputCompute[176]) );
  BUF_X4 U781 ( .A(Row1[177]), .Z(OutputCompute[177]) );
  BUF_X4 U782 ( .A(Row1[178]), .Z(OutputCompute[178]) );
  BUF_X4 U783 ( .A(Row1[179]), .Z(OutputCompute[179]) );
  BUF_X4 U784 ( .A(Row1[180]), .Z(OutputCompute[180]) );
  BUF_X4 U785 ( .A(Row1[181]), .Z(OutputCompute[181]) );
  BUF_X4 U786 ( .A(Row1[182]), .Z(OutputCompute[182]) );
  BUF_X4 U787 ( .A(Row1[183]), .Z(OutputCompute[183]) );
  NAND2_X2 U788 ( .A1(n4800), .A2(n8), .ZN(n51) );
  BUF_X4 U789 ( .A(Row2[248]), .Z(Output_2Row2[248]) );
  BUF_X4 U790 ( .A(Row2[252]), .Z(Output_2Row2[252]) );
  BUF_X4 U791 ( .A(Row2[249]), .Z(Output_2Row2[249]) );
  BUF_X4 U792 ( .A(Row2[250]), .Z(Output_2Row2[250]) );
  BUF_X4 U793 ( .A(Row2[251]), .Z(Output_2Row2[251]) );
  BUF_X4 U794 ( .A(PaddedRow[0]), .Z(WriteBus[0]) );
  BUF_X4 U795 ( .A(Row1[0]), .Z(OutputPaddedRow[0]) );
  BUF_X4 U796 ( .A(PaddedRow[1]), .Z(WriteBus[1]) );
  BUF_X4 U797 ( .A(Row1[1]), .Z(OutputPaddedRow[1]) );
  BUF_X4 U798 ( .A(PaddedRow[2]), .Z(WriteBus[2]) );
  BUF_X4 U799 ( .A(Row1[2]), .Z(OutputPaddedRow[2]) );
  BUF_X4 U800 ( .A(PaddedRow[3]), .Z(WriteBus[3]) );
  BUF_X4 U801 ( .A(Row1[3]), .Z(OutputPaddedRow[3]) );
  BUF_X4 U802 ( .A(PaddedRow[4]), .Z(WriteBus[4]) );
  BUF_X4 U803 ( .A(Row1[4]), .Z(OutputPaddedRow[4]) );
  BUF_X4 U804 ( .A(PaddedRow[5]), .Z(WriteBus[5]) );
  BUF_X4 U805 ( .A(Row1[5]), .Z(OutputPaddedRow[5]) );
  BUF_X4 U806 ( .A(PaddedRow[6]), .Z(WriteBus[6]) );
  BUF_X4 U807 ( .A(Row1[6]), .Z(OutputPaddedRow[6]) );
  BUF_X4 U808 ( .A(PaddedRow[7]), .Z(WriteBus[7]) );
  BUF_X4 U809 ( .A(Row1[7]), .Z(OutputPaddedRow[7]) );
  BUF_X4 U810 ( .A(PaddedRow[8]), .Z(WriteBus[8]) );
  BUF_X4 U811 ( .A(Row1[8]), .Z(OutputPaddedRow[8]) );
  BUF_X4 U812 ( .A(PaddedRow[9]), .Z(WriteBus[9]) );
  BUF_X4 U813 ( .A(Row1[9]), .Z(OutputPaddedRow[9]) );
  BUF_X4 U814 ( .A(PaddedRow[10]), .Z(WriteBus[10]) );
  BUF_X4 U815 ( .A(Row1[10]), .Z(OutputPaddedRow[10]) );
  BUF_X4 U816 ( .A(PaddedRow[11]), .Z(WriteBus[11]) );
  BUF_X4 U817 ( .A(Row1[11]), .Z(OutputPaddedRow[11]) );
  BUF_X4 U818 ( .A(PaddedRow[12]), .Z(WriteBus[12]) );
  BUF_X4 U819 ( .A(Row1[12]), .Z(OutputPaddedRow[12]) );
  BUF_X4 U820 ( .A(PaddedRow[13]), .Z(WriteBus[13]) );
  BUF_X4 U821 ( .A(Row1[13]), .Z(OutputPaddedRow[13]) );
  BUF_X4 U822 ( .A(PaddedRow[14]), .Z(WriteBus[14]) );
  BUF_X4 U823 ( .A(Row1[14]), .Z(OutputPaddedRow[14]) );
  BUF_X4 U824 ( .A(PaddedRow[15]), .Z(WriteBus[15]) );
  BUF_X4 U825 ( .A(Row1[15]), .Z(OutputPaddedRow[15]) );
  BUF_X4 U826 ( .A(PaddedRow[16]), .Z(WriteBus[16]) );
  BUF_X4 U827 ( .A(Row1[16]), .Z(OutputPaddedRow[16]) );
  BUF_X4 U828 ( .A(PaddedRow[17]), .Z(WriteBus[17]) );
  BUF_X4 U829 ( .A(Row1[17]), .Z(OutputPaddedRow[17]) );
  BUF_X4 U830 ( .A(PaddedRow[18]), .Z(WriteBus[18]) );
  BUF_X4 U831 ( .A(Row1[18]), .Z(OutputPaddedRow[18]) );
  BUF_X4 U832 ( .A(PaddedRow[19]), .Z(WriteBus[19]) );
  BUF_X4 U833 ( .A(Row1[19]), .Z(OutputPaddedRow[19]) );
  BUF_X4 U834 ( .A(PaddedRow[20]), .Z(WriteBus[20]) );
  BUF_X4 U835 ( .A(Row1[20]), .Z(OutputPaddedRow[20]) );
  BUF_X4 U836 ( .A(PaddedRow[21]), .Z(WriteBus[21]) );
  BUF_X4 U837 ( .A(Row1[21]), .Z(OutputPaddedRow[21]) );
  BUF_X4 U838 ( .A(PaddedRow[22]), .Z(WriteBus[22]) );
  BUF_X4 U839 ( .A(Row1[22]), .Z(OutputPaddedRow[22]) );
  BUF_X4 U840 ( .A(PaddedRow[23]), .Z(WriteBus[23]) );
  BUF_X4 U841 ( .A(Row1[23]), .Z(OutputPaddedRow[23]) );
  BUF_X4 U842 ( .A(PaddedRow[24]), .Z(WriteBus[24]) );
  BUF_X4 U843 ( .A(Row1[24]), .Z(OutputPaddedRow[24]) );
  BUF_X4 U844 ( .A(PaddedRow[25]), .Z(WriteBus[25]) );
  BUF_X4 U845 ( .A(Row1[25]), .Z(OutputPaddedRow[25]) );
  BUF_X4 U846 ( .A(PaddedRow[26]), .Z(WriteBus[26]) );
  BUF_X4 U847 ( .A(Row1[26]), .Z(OutputPaddedRow[26]) );
  BUF_X4 U848 ( .A(PaddedRow[27]), .Z(WriteBus[27]) );
  BUF_X4 U849 ( .A(Row1[27]), .Z(OutputPaddedRow[27]) );
  BUF_X4 U850 ( .A(PaddedRow[28]), .Z(WriteBus[28]) );
  BUF_X4 U851 ( .A(Row1[28]), .Z(OutputPaddedRow[28]) );
  BUF_X4 U852 ( .A(PaddedRow[29]), .Z(WriteBus[29]) );
  BUF_X4 U853 ( .A(Row1[29]), .Z(OutputPaddedRow[29]) );
  BUF_X4 U854 ( .A(PaddedRow[30]), .Z(WriteBus[30]) );
  BUF_X4 U855 ( .A(Row1[30]), .Z(OutputPaddedRow[30]) );
  BUF_X4 U856 ( .A(PaddedRow[31]), .Z(WriteBus[31]) );
  BUF_X4 U857 ( .A(Row1[31]), .Z(OutputPaddedRow[31]) );
  BUF_X4 U858 ( .A(PaddedRow[32]), .Z(WriteBus[32]) );
  BUF_X4 U859 ( .A(Row1[32]), .Z(OutputPaddedRow[32]) );
  BUF_X4 U860 ( .A(PaddedRow[33]), .Z(WriteBus[33]) );
  BUF_X4 U861 ( .A(Row1[33]), .Z(OutputPaddedRow[33]) );
  BUF_X4 U862 ( .A(PaddedRow[34]), .Z(WriteBus[34]) );
  BUF_X4 U863 ( .A(Row1[34]), .Z(OutputPaddedRow[34]) );
  BUF_X4 U864 ( .A(PaddedRow[35]), .Z(WriteBus[35]) );
  BUF_X4 U865 ( .A(Row1[35]), .Z(OutputPaddedRow[35]) );
  BUF_X4 U866 ( .A(PaddedRow[36]), .Z(WriteBus[36]) );
  BUF_X4 U867 ( .A(Row1[36]), .Z(OutputPaddedRow[36]) );
  BUF_X4 U868 ( .A(PaddedRow[37]), .Z(WriteBus[37]) );
  BUF_X4 U869 ( .A(Row1[37]), .Z(OutputPaddedRow[37]) );
  BUF_X4 U870 ( .A(PaddedRow[38]), .Z(WriteBus[38]) );
  BUF_X4 U871 ( .A(Row1[38]), .Z(OutputPaddedRow[38]) );
  BUF_X4 U872 ( .A(PaddedRow[39]), .Z(WriteBus[39]) );
  BUF_X4 U873 ( .A(Row1[39]), .Z(OutputPaddedRow[39]) );
  BUF_X4 U874 ( .A(PaddedRow[40]), .Z(WriteBus[40]) );
  BUF_X4 U875 ( .A(Row1[40]), .Z(OutputPaddedRow[40]) );
  BUF_X4 U876 ( .A(PaddedRow[41]), .Z(WriteBus[41]) );
  BUF_X4 U877 ( .A(Row1[41]), .Z(OutputPaddedRow[41]) );
  BUF_X4 U878 ( .A(PaddedRow[42]), .Z(WriteBus[42]) );
  BUF_X4 U879 ( .A(Row1[42]), .Z(OutputPaddedRow[42]) );
  BUF_X4 U880 ( .A(PaddedRow[43]), .Z(WriteBus[43]) );
  BUF_X4 U881 ( .A(Row1[43]), .Z(OutputPaddedRow[43]) );
  BUF_X4 U882 ( .A(PaddedRow[44]), .Z(WriteBus[44]) );
  BUF_X4 U883 ( .A(Row1[44]), .Z(OutputPaddedRow[44]) );
  BUF_X4 U884 ( .A(PaddedRow[45]), .Z(WriteBus[45]) );
  BUF_X4 U885 ( .A(Row1[45]), .Z(OutputPaddedRow[45]) );
  BUF_X4 U886 ( .A(PaddedRow[46]), .Z(WriteBus[46]) );
  BUF_X4 U887 ( .A(Row1[46]), .Z(OutputPaddedRow[46]) );
  BUF_X4 U888 ( .A(PaddedRow[47]), .Z(WriteBus[47]) );
  BUF_X4 U889 ( .A(Row1[47]), .Z(OutputPaddedRow[47]) );
  BUF_X4 U890 ( .A(PaddedRow[75]), .Z(WriteBus[75]) );
  BUF_X4 U891 ( .A(Row1[75]), .Z(OutputPaddedRow[75]) );
  BUF_X4 U892 ( .A(PaddedRow[76]), .Z(WriteBus[76]) );
  BUF_X4 U893 ( .A(Row1[76]), .Z(OutputPaddedRow[76]) );
  BUF_X4 U894 ( .A(PaddedRow[77]), .Z(WriteBus[77]) );
  BUF_X4 U895 ( .A(Row1[77]), .Z(OutputPaddedRow[77]) );
  BUF_X4 U896 ( .A(PaddedRow[78]), .Z(WriteBus[78]) );
  BUF_X4 U897 ( .A(Row1[78]), .Z(OutputPaddedRow[78]) );
  BUF_X4 U898 ( .A(PaddedRow[79]), .Z(WriteBus[79]) );
  BUF_X4 U899 ( .A(Row1[79]), .Z(OutputPaddedRow[79]) );
  BUF_X4 U900 ( .A(PaddedRow[107]), .Z(WriteBus[107]) );
  BUF_X4 U901 ( .A(Row1[107]), .Z(OutputPaddedRow[107]) );
  BUF_X4 U902 ( .A(PaddedRow[108]), .Z(WriteBus[108]) );
  BUF_X4 U903 ( .A(Row1[108]), .Z(OutputPaddedRow[108]) );
  BUF_X4 U904 ( .A(PaddedRow[109]), .Z(WriteBus[109]) );
  BUF_X4 U905 ( .A(Row1[109]), .Z(OutputPaddedRow[109]) );
  BUF_X4 U906 ( .A(PaddedRow[110]), .Z(WriteBus[110]) );
  BUF_X4 U907 ( .A(Row1[110]), .Z(OutputPaddedRow[110]) );
  BUF_X4 U908 ( .A(PaddedRow[111]), .Z(WriteBus[111]) );
  BUF_X4 U909 ( .A(Row1[111]), .Z(OutputPaddedRow[111]) );
  BUF_X4 U910 ( .A(PaddedRow[192]), .Z(WriteBus[192]) );
  BUF_X4 U911 ( .A(Row1[192]), .Z(OutputPaddedRow[192]) );
  BUF_X4 U912 ( .A(PaddedRow[193]), .Z(WriteBus[193]) );
  BUF_X4 U913 ( .A(Row1[193]), .Z(OutputPaddedRow[193]) );
  BUF_X4 U914 ( .A(PaddedRow[194]), .Z(WriteBus[194]) );
  BUF_X4 U915 ( .A(Row1[194]), .Z(OutputPaddedRow[194]) );
  BUF_X4 U916 ( .A(PaddedRow[195]), .Z(WriteBus[195]) );
  BUF_X4 U917 ( .A(Row1[195]), .Z(OutputPaddedRow[195]) );
  BUF_X4 U918 ( .A(PaddedRow[196]), .Z(WriteBus[196]) );
  BUF_X4 U919 ( .A(Row1[196]), .Z(OutputPaddedRow[196]) );
  BUF_X4 U920 ( .A(PaddedRow[197]), .Z(WriteBus[197]) );
  BUF_X4 U921 ( .A(Row1[197]), .Z(OutputPaddedRow[197]) );
  BUF_X4 U922 ( .A(PaddedRow[198]), .Z(WriteBus[198]) );
  BUF_X4 U923 ( .A(Row1[198]), .Z(OutputPaddedRow[198]) );
  BUF_X4 U924 ( .A(PaddedRow[199]), .Z(WriteBus[199]) );
  BUF_X4 U925 ( .A(Row1[199]), .Z(OutputPaddedRow[199]) );
  BUF_X4 U926 ( .A(PaddedRow[200]), .Z(WriteBus[200]) );
  BUF_X4 U927 ( .A(Row1[200]), .Z(OutputPaddedRow[200]) );
  BUF_X4 U928 ( .A(PaddedRow[201]), .Z(WriteBus[201]) );
  BUF_X4 U929 ( .A(Row1[201]), .Z(OutputPaddedRow[201]) );
  BUF_X4 U930 ( .A(PaddedRow[202]), .Z(WriteBus[202]) );
  BUF_X4 U931 ( .A(Row1[202]), .Z(OutputPaddedRow[202]) );
  BUF_X4 U932 ( .A(PaddedRow[203]), .Z(WriteBus[203]) );
  BUF_X4 U933 ( .A(Row1[203]), .Z(OutputPaddedRow[203]) );
  BUF_X4 U934 ( .A(PaddedRow[204]), .Z(WriteBus[204]) );
  BUF_X4 U935 ( .A(Row1[204]), .Z(OutputPaddedRow[204]) );
  BUF_X4 U936 ( .A(PaddedRow[205]), .Z(WriteBus[205]) );
  BUF_X4 U937 ( .A(Row1[205]), .Z(OutputPaddedRow[205]) );
  BUF_X4 U938 ( .A(PaddedRow[206]), .Z(WriteBus[206]) );
  BUF_X4 U939 ( .A(Row1[206]), .Z(OutputPaddedRow[206]) );
  BUF_X4 U940 ( .A(PaddedRow[207]), .Z(WriteBus[207]) );
  BUF_X4 U941 ( .A(Row1[207]), .Z(OutputPaddedRow[207]) );
  BUF_X4 U942 ( .A(PaddedRow[208]), .Z(WriteBus[208]) );
  BUF_X4 U943 ( .A(Row1[208]), .Z(OutputPaddedRow[208]) );
  BUF_X4 U944 ( .A(PaddedRow[209]), .Z(WriteBus[209]) );
  BUF_X4 U945 ( .A(Row1[209]), .Z(OutputPaddedRow[209]) );
  BUF_X4 U946 ( .A(PaddedRow[210]), .Z(WriteBus[210]) );
  BUF_X4 U947 ( .A(Row1[210]), .Z(OutputPaddedRow[210]) );
  BUF_X4 U948 ( .A(PaddedRow[211]), .Z(WriteBus[211]) );
  BUF_X4 U949 ( .A(Row1[211]), .Z(OutputPaddedRow[211]) );
  BUF_X4 U950 ( .A(PaddedRow[212]), .Z(WriteBus[212]) );
  BUF_X4 U951 ( .A(Row1[212]), .Z(OutputPaddedRow[212]) );
  BUF_X4 U952 ( .A(PaddedRow[213]), .Z(WriteBus[213]) );
  BUF_X4 U953 ( .A(Row1[213]), .Z(OutputPaddedRow[213]) );
  BUF_X4 U954 ( .A(PaddedRow[214]), .Z(WriteBus[214]) );
  BUF_X4 U955 ( .A(Row1[214]), .Z(OutputPaddedRow[214]) );
  BUF_X4 U956 ( .A(PaddedRow[215]), .Z(WriteBus[215]) );
  BUF_X4 U957 ( .A(Row1[215]), .Z(OutputPaddedRow[215]) );
  BUF_X4 U958 ( .A(PaddedRow[216]), .Z(WriteBus[216]) );
  BUF_X4 U959 ( .A(Row1[216]), .Z(OutputPaddedRow[216]) );
  BUF_X4 U960 ( .A(PaddedRow[217]), .Z(WriteBus[217]) );
  BUF_X4 U961 ( .A(Row1[217]), .Z(OutputPaddedRow[217]) );
  BUF_X4 U962 ( .A(PaddedRow[218]), .Z(WriteBus[218]) );
  BUF_X4 U963 ( .A(Row1[218]), .Z(OutputPaddedRow[218]) );
  BUF_X4 U964 ( .A(PaddedRow[219]), .Z(WriteBus[219]) );
  BUF_X4 U965 ( .A(Row1[219]), .Z(OutputPaddedRow[219]) );
  BUF_X4 U966 ( .A(PaddedRow[220]), .Z(WriteBus[220]) );
  BUF_X4 U967 ( .A(Row1[220]), .Z(OutputPaddedRow[220]) );
  BUF_X4 U968 ( .A(PaddedRow[221]), .Z(WriteBus[221]) );
  BUF_X4 U969 ( .A(Row1[221]), .Z(OutputPaddedRow[221]) );
  BUF_X4 U970 ( .A(PaddedRow[222]), .Z(WriteBus[222]) );
  BUF_X4 U971 ( .A(Row1[222]), .Z(OutputPaddedRow[222]) );
  BUF_X4 U972 ( .A(PaddedRow[223]), .Z(WriteBus[223]) );
  BUF_X4 U973 ( .A(Row1[223]), .Z(OutputPaddedRow[223]) );
  BUF_X4 U974 ( .A(PaddedRow[224]), .Z(WriteBus[224]) );
  BUF_X4 U975 ( .A(Row1[224]), .Z(OutputPaddedRow[224]) );
  BUF_X4 U976 ( .A(PaddedRow[225]), .Z(WriteBus[225]) );
  BUF_X4 U977 ( .A(Row1[225]), .Z(OutputPaddedRow[225]) );
  BUF_X4 U978 ( .A(PaddedRow[226]), .Z(WriteBus[226]) );
  BUF_X4 U979 ( .A(Row1[226]), .Z(OutputPaddedRow[226]) );
  BUF_X4 U980 ( .A(PaddedRow[227]), .Z(WriteBus[227]) );
  BUF_X4 U981 ( .A(Row1[227]), .Z(OutputPaddedRow[227]) );
  BUF_X4 U982 ( .A(PaddedRow[228]), .Z(WriteBus[228]) );
  BUF_X4 U983 ( .A(Row1[228]), .Z(OutputPaddedRow[228]) );
  BUF_X4 U984 ( .A(PaddedRow[229]), .Z(WriteBus[229]) );
  BUF_X4 U985 ( .A(Row1[229]), .Z(OutputPaddedRow[229]) );
  BUF_X4 U986 ( .A(PaddedRow[230]), .Z(WriteBus[230]) );
  BUF_X4 U987 ( .A(Row1[230]), .Z(OutputPaddedRow[230]) );
  BUF_X4 U988 ( .A(PaddedRow[231]), .Z(WriteBus[231]) );
  BUF_X4 U989 ( .A(Row1[231]), .Z(OutputPaddedRow[231]) );
  BUF_X4 U990 ( .A(PaddedRow[232]), .Z(WriteBus[232]) );
  BUF_X4 U991 ( .A(Row1[232]), .Z(OutputPaddedRow[232]) );
  BUF_X4 U992 ( .A(PaddedRow[233]), .Z(WriteBus[233]) );
  BUF_X4 U993 ( .A(Row1[233]), .Z(OutputPaddedRow[233]) );
  BUF_X4 U994 ( .A(PaddedRow[234]), .Z(WriteBus[234]) );
  BUF_X4 U995 ( .A(Row1[234]), .Z(OutputPaddedRow[234]) );
  BUF_X4 U996 ( .A(PaddedRow[235]), .Z(WriteBus[235]) );
  BUF_X4 U997 ( .A(Row1[235]), .Z(OutputPaddedRow[235]) );
  BUF_X4 U998 ( .A(PaddedRow[236]), .Z(WriteBus[236]) );
  BUF_X4 U999 ( .A(Row1[236]), .Z(OutputPaddedRow[236]) );
  BUF_X4 U1000 ( .A(PaddedRow[237]), .Z(WriteBus[237]) );
  BUF_X4 U1001 ( .A(Row1[237]), .Z(OutputPaddedRow[237]) );
  BUF_X4 U1002 ( .A(PaddedRow[238]), .Z(WriteBus[238]) );
  BUF_X4 U1003 ( .A(Row1[238]), .Z(OutputPaddedRow[238]) );
  BUF_X4 U1004 ( .A(PaddedRow[239]), .Z(WriteBus[239]) );
  BUF_X4 U1005 ( .A(Row1[239]), .Z(OutputPaddedRow[239]) );
  BUF_X4 U1006 ( .A(Row1[111]), .Z(Output_2Row1[111]) );
  BUF_X4 U1007 ( .A(Row1[75]), .Z(Output_2Row1[75]) );
  BUF_X4 U1008 ( .A(Row1[76]), .Z(Output_2Row1[76]) );
  BUF_X4 U1009 ( .A(Row1[77]), .Z(Output_2Row1[77]) );
  BUF_X4 U1010 ( .A(Row1[78]), .Z(Output_2Row1[78]) );
  BUF_X4 U1011 ( .A(Row1[79]), .Z(Output_2Row1[79]) );
  BUF_X4 U1012 ( .A(Row1[91]), .Z(Output_2Row1[91]) );
  BUF_X4 U1013 ( .A(Row1[92]), .Z(Output_2Row1[92]) );
  BUF_X4 U1014 ( .A(Row1[93]), .Z(Output_2Row1[93]) );
  BUF_X4 U1015 ( .A(Row1[94]), .Z(Output_2Row1[94]) );
  BUF_X4 U1016 ( .A(Row1[95]), .Z(Output_2Row1[95]) );
  BUF_X4 U1017 ( .A(Row1[107]), .Z(Output_2Row1[107]) );
  BUF_X4 U1018 ( .A(Row1[108]), .Z(Output_2Row1[108]) );
  BUF_X4 U1019 ( .A(Row1[109]), .Z(Output_2Row1[109]) );
  BUF_X4 U1020 ( .A(Row1[110]), .Z(Output_2Row1[110]) );
  BUF_X4 U1021 ( .A(Row1[0]), .Z(Output_2Row1[0]) );
  BUF_X4 U1022 ( .A(Row1[1]), .Z(Output_2Row1[1]) );
  BUF_X4 U1023 ( .A(Row1[2]), .Z(Output_2Row1[2]) );
  BUF_X4 U1024 ( .A(Row1[3]), .Z(Output_2Row1[3]) );
  BUF_X4 U1025 ( .A(Row1[4]), .Z(Output_2Row1[4]) );
  BUF_X4 U1026 ( .A(Row1[5]), .Z(Output_2Row1[5]) );
  BUF_X4 U1027 ( .A(Row1[6]), .Z(Output_2Row1[6]) );
  BUF_X4 U1028 ( .A(Row1[7]), .Z(Output_2Row1[7]) );
  BUF_X4 U1029 ( .A(Row1[8]), .Z(Output_2Row1[8]) );
  BUF_X4 U1030 ( .A(Row1[9]), .Z(Output_2Row1[9]) );
  BUF_X4 U1031 ( .A(Row1[10]), .Z(Output_2Row1[10]) );
  BUF_X4 U1032 ( .A(Row1[11]), .Z(Output_2Row1[11]) );
  BUF_X4 U1033 ( .A(Row1[12]), .Z(Output_2Row1[12]) );
  BUF_X4 U1034 ( .A(Row1[13]), .Z(Output_2Row1[13]) );
  BUF_X4 U1035 ( .A(Row1[14]), .Z(Output_2Row1[14]) );
  BUF_X4 U1036 ( .A(Row1[15]), .Z(Output_2Row1[15]) );
  BUF_X4 U1037 ( .A(Row1[16]), .Z(Output_2Row1[16]) );
  BUF_X4 U1038 ( .A(Row1[17]), .Z(Output_2Row1[17]) );
  BUF_X4 U1039 ( .A(Row1[18]), .Z(Output_2Row1[18]) );
  BUF_X4 U1040 ( .A(Row1[19]), .Z(Output_2Row1[19]) );
  BUF_X4 U1041 ( .A(Row1[20]), .Z(Output_2Row1[20]) );
  BUF_X4 U1042 ( .A(Row1[21]), .Z(Output_2Row1[21]) );
  BUF_X4 U1043 ( .A(Row1[22]), .Z(Output_2Row1[22]) );
  BUF_X4 U1044 ( .A(Row1[23]), .Z(Output_2Row1[23]) );
  BUF_X4 U1045 ( .A(Row1[24]), .Z(Output_2Row1[24]) );
  BUF_X4 U1046 ( .A(Row1[25]), .Z(Output_2Row1[25]) );
  BUF_X4 U1047 ( .A(Row1[26]), .Z(Output_2Row1[26]) );
  BUF_X4 U1048 ( .A(Row1[27]), .Z(Output_2Row1[27]) );
  BUF_X4 U1049 ( .A(Row1[28]), .Z(Output_2Row1[28]) );
  BUF_X4 U1050 ( .A(Row1[29]), .Z(Output_2Row1[29]) );
  BUF_X4 U1051 ( .A(Row1[30]), .Z(Output_2Row1[30]) );
  BUF_X4 U1052 ( .A(Row1[31]), .Z(Output_2Row1[31]) );
  BUF_X4 U1053 ( .A(Row1[32]), .Z(Output_2Row1[32]) );
  BUF_X4 U1054 ( .A(Row1[33]), .Z(Output_2Row1[33]) );
  BUF_X4 U1055 ( .A(Row1[34]), .Z(Output_2Row1[34]) );
  BUF_X4 U1056 ( .A(Row1[35]), .Z(Output_2Row1[35]) );
  BUF_X4 U1057 ( .A(Row1[36]), .Z(Output_2Row1[36]) );
  BUF_X4 U1058 ( .A(Row1[37]), .Z(Output_2Row1[37]) );
  BUF_X4 U1059 ( .A(Row1[38]), .Z(Output_2Row1[38]) );
  BUF_X4 U1060 ( .A(Row1[39]), .Z(Output_2Row1[39]) );
  BUF_X4 U1061 ( .A(Row1[40]), .Z(Output_2Row1[40]) );
  BUF_X4 U1062 ( .A(Row1[41]), .Z(Output_2Row1[41]) );
  BUF_X4 U1063 ( .A(Row1[42]), .Z(Output_2Row1[42]) );
  BUF_X4 U1064 ( .A(Row1[43]), .Z(Output_2Row1[43]) );
  BUF_X4 U1065 ( .A(Row1[44]), .Z(Output_2Row1[44]) );
  BUF_X4 U1066 ( .A(Row1[45]), .Z(Output_2Row1[45]) );
  BUF_X4 U1067 ( .A(Row1[46]), .Z(Output_2Row1[46]) );
  BUF_X4 U1068 ( .A(Row1[47]), .Z(Output_2Row1[47]) );
  BUF_X4 U1069 ( .A(Row1[175]), .Z(Output_2Row1[175]) );
  BUF_X4 U1070 ( .A(Row1[128]), .Z(Output_2Row1[128]) );
  BUF_X4 U1071 ( .A(Row1[129]), .Z(Output_2Row1[129]) );
  BUF_X4 U1072 ( .A(Row1[130]), .Z(Output_2Row1[130]) );
  BUF_X4 U1073 ( .A(Row1[131]), .Z(Output_2Row1[131]) );
  BUF_X4 U1074 ( .A(Row1[132]), .Z(Output_2Row1[132]) );
  BUF_X4 U1075 ( .A(Row1[133]), .Z(Output_2Row1[133]) );
  BUF_X4 U1076 ( .A(Row1[134]), .Z(Output_2Row1[134]) );
  BUF_X4 U1077 ( .A(Row1[135]), .Z(Output_2Row1[135]) );
  BUF_X4 U1078 ( .A(Row1[136]), .Z(Output_2Row1[136]) );
  BUF_X4 U1079 ( .A(Row1[137]), .Z(Output_2Row1[137]) );
  BUF_X4 U1080 ( .A(Row1[138]), .Z(Output_2Row1[138]) );
  BUF_X4 U1081 ( .A(Row1[139]), .Z(Output_2Row1[139]) );
  BUF_X4 U1082 ( .A(Row1[140]), .Z(Output_2Row1[140]) );
  BUF_X4 U1083 ( .A(Row1[141]), .Z(Output_2Row1[141]) );
  BUF_X4 U1084 ( .A(Row1[142]), .Z(Output_2Row1[142]) );
  BUF_X4 U1085 ( .A(Row1[143]), .Z(Output_2Row1[143]) );
  BUF_X4 U1086 ( .A(Row1[144]), .Z(Output_2Row1[144]) );
  BUF_X4 U1087 ( .A(Row1[145]), .Z(Output_2Row1[145]) );
  BUF_X4 U1088 ( .A(Row1[146]), .Z(Output_2Row1[146]) );
  BUF_X4 U1089 ( .A(Row1[147]), .Z(Output_2Row1[147]) );
  BUF_X4 U1090 ( .A(Row1[148]), .Z(Output_2Row1[148]) );
  BUF_X4 U1091 ( .A(Row1[149]), .Z(Output_2Row1[149]) );
  BUF_X4 U1092 ( .A(Row1[150]), .Z(Output_2Row1[150]) );
  BUF_X4 U1093 ( .A(Row1[151]), .Z(Output_2Row1[151]) );
  BUF_X4 U1094 ( .A(Row1[152]), .Z(Output_2Row1[152]) );
  BUF_X4 U1095 ( .A(Row1[153]), .Z(Output_2Row1[153]) );
  BUF_X4 U1096 ( .A(Row1[154]), .Z(Output_2Row1[154]) );
  BUF_X4 U1097 ( .A(Row1[155]), .Z(Output_2Row1[155]) );
  BUF_X4 U1098 ( .A(Row1[156]), .Z(Output_2Row1[156]) );
  BUF_X4 U1099 ( .A(Row1[157]), .Z(Output_2Row1[157]) );
  BUF_X4 U1100 ( .A(Row1[158]), .Z(Output_2Row1[158]) );
  BUF_X4 U1101 ( .A(Row1[159]), .Z(Output_2Row1[159]) );
  BUF_X4 U1102 ( .A(Row1[160]), .Z(Output_2Row1[160]) );
  BUF_X4 U1103 ( .A(Row1[161]), .Z(Output_2Row1[161]) );
  BUF_X4 U1104 ( .A(Row1[162]), .Z(Output_2Row1[162]) );
  BUF_X4 U1105 ( .A(Row1[163]), .Z(Output_2Row1[163]) );
  BUF_X4 U1106 ( .A(Row1[164]), .Z(Output_2Row1[164]) );
  BUF_X4 U1107 ( .A(Row1[165]), .Z(Output_2Row1[165]) );
  BUF_X4 U1108 ( .A(Row1[166]), .Z(Output_2Row1[166]) );
  BUF_X4 U1109 ( .A(Row1[167]), .Z(Output_2Row1[167]) );
  BUF_X4 U1110 ( .A(Row1[168]), .Z(Output_2Row1[168]) );
  BUF_X4 U1111 ( .A(Row1[169]), .Z(Output_2Row1[169]) );
  BUF_X4 U1112 ( .A(Row1[170]), .Z(Output_2Row1[170]) );
  BUF_X4 U1113 ( .A(Row1[171]), .Z(Output_2Row1[171]) );
  BUF_X4 U1114 ( .A(Row1[172]), .Z(Output_2Row1[172]) );
  BUF_X4 U1115 ( .A(Row1[173]), .Z(Output_2Row1[173]) );
  BUF_X4 U1116 ( .A(Row1[174]), .Z(Output_2Row1[174]) );
  BUF_X4 U1117 ( .A(Row1[239]), .Z(Output_2Row1[239]) );
  BUF_X4 U1118 ( .A(Row2[246]), .Z(Output_2Row2[246]) );
  BUF_X4 U1119 ( .A(Row2[247]), .Z(Output_2Row2[247]) );
  BUF_X4 U1120 ( .A(Row2[243]), .Z(Output_2Row2[243]) );
  BUF_X4 U1121 ( .A(Row2[240]), .Z(Output_2Row2[240]) );
  BUF_X4 U1122 ( .A(Row2[245]), .Z(Output_2Row2[245]) );
  BUF_X4 U1123 ( .A(Row2[244]), .Z(Output_2Row2[244]) );
  BUF_X4 U1124 ( .A(Row2[242]), .Z(Output_2Row2[242]) );
  BUF_X4 U1125 ( .A(Row2[241]), .Z(Output_2Row2[241]) );
  BUF_X4 U1126 ( .A(Row2[254]), .Z(Output_2Row2[254]) );
  BUF_X4 U1127 ( .A(Row2[253]), .Z(Output_2Row2[253]) );
  BUF_X4 U1128 ( .A(Row2[255]), .Z(Output_2Row2[255]) );
  BUF_X4 U1129 ( .A(PaddedRow[91]), .Z(WriteBus[91]) );
  BUF_X4 U1130 ( .A(Row1[91]), .Z(OutputPaddedRow[91]) );
  BUF_X4 U1131 ( .A(PaddedRow[92]), .Z(WriteBus[92]) );
  BUF_X4 U1132 ( .A(Row1[92]), .Z(OutputPaddedRow[92]) );
  BUF_X4 U1133 ( .A(PaddedRow[93]), .Z(WriteBus[93]) );
  BUF_X4 U1134 ( .A(Row1[93]), .Z(OutputPaddedRow[93]) );
  BUF_X4 U1135 ( .A(PaddedRow[94]), .Z(WriteBus[94]) );
  BUF_X4 U1136 ( .A(Row1[94]), .Z(OutputPaddedRow[94]) );
  BUF_X4 U1137 ( .A(PaddedRow[95]), .Z(WriteBus[95]) );
  BUF_X4 U1138 ( .A(Row1[95]), .Z(OutputPaddedRow[95]) );
  INV_X4 U1139 ( .A(n4770), .ZN(n4769) );
  AOI22_X2 U1140 ( .A1(n83), .A2(\U3/U7/DATA6_0 ), .B1(n84), .B2(
        \U3/U7/DATA5_0 ), .ZN(n114) );
  AOI22_X2 U1141 ( .A1(n85), .A2(\U3/U7/DATA4_0 ), .B1(\U3/U7/DATA3_0 ), .B2(
        n4801), .ZN(n113) );
  AOI222_X1 U1142 ( .A1(\U3/U7/DATA7_0 ), .A2(n1830), .B1(\U3/U7/DATA2_0 ), 
        .B2(n81), .C1(\U3/U7/DATA1_0 ), .C2(n82), .ZN(n115) );
  AOI22_X2 U1143 ( .A1(n83), .A2(\U3/U7/DATA6_1 ), .B1(n84), .B2(
        \U3/U7/DATA5_1 ), .ZN(n111) );
  AOI22_X2 U1144 ( .A1(n85), .A2(\U3/U7/DATA4_1 ), .B1(\U3/U7/DATA3_1 ), .B2(
        n4801), .ZN(n110) );
  AOI222_X1 U1145 ( .A1(\U3/U7/DATA7_1 ), .A2(n1830), .B1(\U3/U7/DATA2_1 ), 
        .B2(n81), .C1(\U3/U7/DATA1_1 ), .C2(n82), .ZN(n112) );
  AOI22_X2 U1146 ( .A1(n83), .A2(\U3/U7/DATA6_2 ), .B1(n84), .B2(
        \U3/U7/DATA5_2 ), .ZN(n105) );
  AOI22_X2 U1147 ( .A1(n85), .A2(\U3/U7/DATA4_2 ), .B1(\U3/U7/DATA3_2 ), .B2(
        n4801), .ZN(n104) );
  AOI222_X1 U1148 ( .A1(\U3/U7/DATA7_2 ), .A2(n1830), .B1(\U3/U7/DATA2_2 ), 
        .B2(n81), .C1(\U3/U7/DATA1_2 ), .C2(n82), .ZN(n106) );
  AOI22_X2 U1149 ( .A1(n83), .A2(\U3/U7/DATA6_3 ), .B1(n84), .B2(
        \U3/U7/DATA5_3 ), .ZN(n102) );
  AOI22_X2 U1150 ( .A1(n85), .A2(\U3/U7/DATA4_3 ), .B1(\U3/U7/DATA3_3 ), .B2(
        n4801), .ZN(n101) );
  AOI222_X1 U1151 ( .A1(\U3/U7/DATA7_3 ), .A2(n1830), .B1(\U3/U7/DATA2_3 ), 
        .B2(n81), .C1(\U3/U7/DATA1_3 ), .C2(n82), .ZN(n103) );
  AOI22_X2 U1152 ( .A1(n83), .A2(\U3/U7/DATA6_4 ), .B1(n84), .B2(
        \U3/U7/DATA5_4 ), .ZN(n99) );
  AOI22_X2 U1153 ( .A1(n85), .A2(\U3/U7/DATA4_4 ), .B1(\U3/U7/DATA3_4 ), .B2(
        n4801), .ZN(n98) );
  AOI222_X1 U1154 ( .A1(\U3/U7/DATA7_4 ), .A2(n1830), .B1(\U3/U7/DATA2_4 ), 
        .B2(n81), .C1(\U3/U7/DATA1_4 ), .C2(n82), .ZN(n100) );
  AOI22_X2 U1155 ( .A1(n83), .A2(\U3/U7/DATA6_5 ), .B1(n84), .B2(
        \U3/U7/DATA5_5 ), .ZN(n96) );
  AOI22_X2 U1156 ( .A1(n85), .A2(\U3/U7/DATA4_5 ), .B1(\U3/U7/DATA3_5 ), .B2(
        n4801), .ZN(n95) );
  AOI222_X1 U1157 ( .A1(\U3/U7/DATA7_5 ), .A2(n1830), .B1(\U3/U7/DATA2_5 ), 
        .B2(n81), .C1(\U3/U7/DATA1_5 ), .C2(n82), .ZN(n97) );
  AOI22_X2 U1158 ( .A1(n83), .A2(\U3/U7/DATA6_6 ), .B1(n84), .B2(
        \U3/U7/DATA5_6 ), .ZN(n93) );
  AOI22_X2 U1159 ( .A1(n85), .A2(\U3/U7/DATA4_6 ), .B1(\U3/U7/DATA3_6 ), .B2(
        n4801), .ZN(n92) );
  AOI222_X1 U1160 ( .A1(\U3/U7/DATA7_6 ), .A2(n1830), .B1(\U3/U7/DATA2_6 ), 
        .B2(n81), .C1(\U3/U7/DATA1_6 ), .C2(n82), .ZN(n94) );
  AOI22_X2 U1161 ( .A1(n83), .A2(\U3/U7/DATA6_7 ), .B1(n84), .B2(
        \U3/U7/DATA5_7 ), .ZN(n90) );
  AOI22_X2 U1162 ( .A1(n85), .A2(\U3/U7/DATA4_7 ), .B1(\U3/U7/DATA3_7 ), .B2(
        n4801), .ZN(n89) );
  AOI222_X1 U1163 ( .A1(\U3/U7/DATA7_7 ), .A2(n1830), .B1(\U3/U7/DATA2_7 ), 
        .B2(n81), .C1(\U3/U7/DATA1_7 ), .C2(n82), .ZN(n91) );
  AOI22_X2 U1164 ( .A1(n83), .A2(\U3/U7/DATA6_8 ), .B1(n84), .B2(
        \U3/U7/DATA5_8 ), .ZN(n87) );
  AOI22_X2 U1165 ( .A1(n85), .A2(\U3/U7/DATA4_8 ), .B1(\U3/U7/DATA3_8 ), .B2(
        n4801), .ZN(n86) );
  AOI222_X1 U1166 ( .A1(\U3/U7/DATA7_8 ), .A2(n1830), .B1(\U3/U7/DATA2_8 ), 
        .B2(n81), .C1(\U3/U7/DATA1_8 ), .C2(n82), .ZN(n88) );
  AOI22_X2 U1167 ( .A1(n83), .A2(\U3/U7/DATA6_9 ), .B1(n84), .B2(
        \U3/U7/DATA5_9 ), .ZN(n79) );
  AOI22_X2 U1168 ( .A1(n85), .A2(\U3/U7/DATA4_9 ), .B1(\U3/U7/DATA3_9 ), .B2(
        n4801), .ZN(n78) );
  AOI222_X1 U1169 ( .A1(\U3/U7/DATA7_9 ), .A2(n1830), .B1(\U3/U7/DATA2_9 ), 
        .B2(n81), .C1(\U3/U7/DATA1_9 ), .C2(n82), .ZN(n80) );
  AOI22_X2 U1170 ( .A1(n83), .A2(\U3/U7/DATA6_10 ), .B1(n84), .B2(
        \U3/U7/DATA5_10 ), .ZN(n108) );
  AOI22_X2 U1171 ( .A1(n85), .A2(\U3/U7/DATA4_10 ), .B1(\U3/U7/DATA3_10 ), 
        .B2(n4801), .ZN(n107) );
  AOI222_X1 U1172 ( .A1(\U3/U7/DATA7_10 ), .A2(n1830), .B1(\U3/U7/DATA2_10 ), 
        .B2(n81), .C1(\U3/U7/DATA1_10 ), .C2(n82), .ZN(n109) );
  AOI222_X1 U1173 ( .A1(\U3/U5/DATA1_2 ), .A2(n2959), .B1(\U3/U5/DATA2_2 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_2 ), .C2(n2958), .ZN(n152) );
  AOI222_X1 U1174 ( .A1(\U3/U5/DATA1_3 ), .A2(n2959), .B1(\U3/U5/DATA2_3 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_3 ), .C2(n2958), .ZN(n141) );
  AOI222_X1 U1175 ( .A1(\U3/U5/DATA1_20 ), .A2(n2959), .B1(\U3/U5/DATA2_20 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_20 ), .C2(n2958), .ZN(n151) );
  AOI222_X1 U1176 ( .A1(\U3/U5/DATA1_21 ), .A2(n2959), .B1(\U3/U5/DATA2_21 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_21 ), .C2(n2958), .ZN(n150) );
  AOI222_X1 U1177 ( .A1(\U3/U5/DATA1_22 ), .A2(n2959), .B1(\U3/U5/DATA2_22 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_22 ), .C2(n2958), .ZN(n149) );
  AOI222_X1 U1178 ( .A1(\U3/U5/DATA1_23 ), .A2(n2959), .B1(\U3/U5/DATA2_23 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_23 ), .C2(n2958), .ZN(n148) );
  AOI222_X1 U1179 ( .A1(\U3/U5/DATA1_24 ), .A2(n2959), .B1(\U3/U5/DATA2_24 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_24 ), .C2(n2958), .ZN(n147) );
  AOI222_X1 U1180 ( .A1(\U3/U5/DATA1_25 ), .A2(n2959), .B1(\U3/U5/DATA2_25 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_25 ), .C2(n2958), .ZN(n146) );
  AOI222_X1 U1181 ( .A1(\U3/U5/DATA1_26 ), .A2(n2959), .B1(\U3/U5/DATA2_26 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_26 ), .C2(n2958), .ZN(n145) );
  AOI222_X1 U1182 ( .A1(\U3/U5/DATA1_27 ), .A2(n2959), .B1(\U3/U5/DATA2_27 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_27 ), .C2(n2958), .ZN(n144) );
  AOI222_X1 U1183 ( .A1(\U3/U5/DATA1_28 ), .A2(n2959), .B1(\U3/U5/DATA2_28 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_28 ), .C2(n2958), .ZN(n143) );
  AOI222_X1 U1184 ( .A1(\U3/U5/DATA1_29 ), .A2(n2959), .B1(\U3/U5/DATA2_29 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_29 ), .C2(n2958), .ZN(n142) );
  BUF_X4 U1185 ( .A(Row2[224]), .Z(Output_1Row2[224]) );
  BUF_X4 U1186 ( .A(Row2[240]), .Z(Output_1Row2[240]) );
  BUF_X4 U1187 ( .A(Row2[96]), .Z(Output_1Row2[96]) );
  BUF_X4 U1188 ( .A(Row2[112]), .Z(Output_1Row2[112]) );
  BUF_X4 U1189 ( .A(Row1[224]), .Z(Output_1Row1[224]) );
  BUF_X4 U1190 ( .A(Row1[240]), .Z(Output_1Row1[240]) );
  BUF_X4 U1191 ( .A(Row2[192]), .Z(Output_1Row2[192]) );
  BUF_X4 U1192 ( .A(Row2[208]), .Z(Output_1Row2[208]) );
  BUF_X4 U1193 ( .A(Row2[64]), .Z(Output_1Row2[64]) );
  BUF_X4 U1194 ( .A(Row2[80]), .Z(Output_1Row2[80]) );
  BUF_X4 U1195 ( .A(Row1[192]), .Z(Output_1Row1[192]) );
  BUF_X4 U1196 ( .A(Row1[208]), .Z(Output_1Row1[208]) );
  BUF_X4 U1197 ( .A(Row2[128]), .Z(Output_1Row2[128]) );
  BUF_X4 U1198 ( .A(Row2[144]), .Z(Output_1Row2[144]) );
  BUF_X4 U1199 ( .A(Row2[0]), .Z(Output_1Row2[0]) );
  BUF_X4 U1200 ( .A(Row2[16]), .Z(Output_1Row2[16]) );
  BUF_X4 U1201 ( .A(Row1[128]), .Z(Output_1Row1[128]) );
  BUF_X4 U1202 ( .A(Row1[144]), .Z(Output_1Row1[144]) );
  BUF_X4 U1203 ( .A(Row1[0]), .Z(Output_1Row1[0]) );
  BUF_X4 U1204 ( .A(Row1[16]), .Z(Output_1Row1[16]) );
  BUF_X4 U1205 ( .A(Row2[170]), .Z(Output_1Row2[170]) );
  BUF_X4 U1206 ( .A(Row2[186]), .Z(Output_1Row2[186]) );
  BUF_X4 U1207 ( .A(Row2[42]), .Z(Output_1Row2[42]) );
  BUF_X4 U1208 ( .A(Row2[58]), .Z(Output_1Row2[58]) );
  BUF_X4 U1209 ( .A(Row2[160]), .Z(Output_1Row2[160]) );
  BUF_X4 U1210 ( .A(Row2[176]), .Z(Output_1Row2[176]) );
  BUF_X4 U1211 ( .A(Row2[32]), .Z(Output_1Row2[32]) );
  BUF_X4 U1212 ( .A(Row2[48]), .Z(Output_1Row2[48]) );
  BUF_X4 U1213 ( .A(Row1[170]), .Z(Output_1Row1[170]) );
  BUF_X4 U1214 ( .A(Row1[186]), .Z(Output_1Row1[186]) );
  BUF_X4 U1215 ( .A(Row1[42]), .Z(Output_1Row1[42]) );
  BUF_X4 U1216 ( .A(Row1[58]), .Z(Output_1Row1[58]) );
  BUF_X4 U1217 ( .A(Row1[160]), .Z(Output_1Row1[160]) );
  BUF_X4 U1218 ( .A(Row1[176]), .Z(Output_1Row1[176]) );
  BUF_X4 U1219 ( .A(Row1[32]), .Z(Output_1Row1[32]) );
  BUF_X4 U1220 ( .A(Row1[48]), .Z(Output_1Row1[48]) );
  OAI21_X2 U1221 ( .B1(n1828), .B2(EOC_Flag), .A(n51), .ZN(n50) );
  BUF_X4 U1222 ( .A(Row2[73]), .Z(Output_1Row2[73]) );
  BUF_X4 U1223 ( .A(Row2[89]), .Z(Output_1Row2[89]) );
  BUF_X4 U1224 ( .A(Row2[72]), .Z(Output_1Row2[72]) );
  BUF_X4 U1225 ( .A(Row2[88]), .Z(Output_1Row2[88]) );
  BUF_X4 U1226 ( .A(Row2[71]), .Z(Output_1Row2[71]) );
  BUF_X4 U1227 ( .A(Row2[87]), .Z(Output_1Row2[87]) );
  BUF_X4 U1228 ( .A(Row2[70]), .Z(Output_1Row2[70]) );
  BUF_X4 U1229 ( .A(Row2[86]), .Z(Output_1Row2[86]) );
  BUF_X4 U1230 ( .A(Row2[69]), .Z(Output_1Row2[69]) );
  BUF_X4 U1231 ( .A(Row2[85]), .Z(Output_1Row2[85]) );
  BUF_X4 U1232 ( .A(Row2[68]), .Z(Output_1Row2[68]) );
  BUF_X4 U1233 ( .A(Row2[84]), .Z(Output_1Row2[84]) );
  BUF_X4 U1234 ( .A(Row2[67]), .Z(Output_1Row2[67]) );
  BUF_X4 U1235 ( .A(Row2[83]), .Z(Output_1Row2[83]) );
  BUF_X4 U1236 ( .A(Row2[66]), .Z(Output_1Row2[66]) );
  BUF_X4 U1237 ( .A(Row2[82]), .Z(Output_1Row2[82]) );
  BUF_X4 U1238 ( .A(Row2[65]), .Z(Output_1Row2[65]) );
  BUF_X4 U1239 ( .A(Row2[81]), .Z(Output_1Row2[81]) );
  BUF_X4 U1240 ( .A(Row2[105]), .Z(Output_1Row2[105]) );
  BUF_X4 U1241 ( .A(Row2[121]), .Z(Output_1Row2[121]) );
  BUF_X4 U1242 ( .A(Row2[104]), .Z(Output_1Row2[104]) );
  BUF_X4 U1243 ( .A(Row2[120]), .Z(Output_1Row2[120]) );
  BUF_X4 U1244 ( .A(Row2[103]), .Z(Output_1Row2[103]) );
  BUF_X4 U1245 ( .A(Row2[119]), .Z(Output_1Row2[119]) );
  BUF_X4 U1246 ( .A(Row2[102]), .Z(Output_1Row2[102]) );
  BUF_X4 U1247 ( .A(Row2[118]), .Z(Output_1Row2[118]) );
  BUF_X4 U1248 ( .A(Row2[101]), .Z(Output_1Row2[101]) );
  BUF_X4 U1249 ( .A(Row2[117]), .Z(Output_1Row2[117]) );
  BUF_X4 U1250 ( .A(Row2[100]), .Z(Output_1Row2[100]) );
  BUF_X4 U1251 ( .A(Row2[116]), .Z(Output_1Row2[116]) );
  BUF_X4 U1252 ( .A(Row2[99]), .Z(Output_1Row2[99]) );
  BUF_X4 U1253 ( .A(Row2[115]), .Z(Output_1Row2[115]) );
  BUF_X4 U1254 ( .A(Row2[98]), .Z(Output_1Row2[98]) );
  BUF_X4 U1255 ( .A(Row2[114]), .Z(Output_1Row2[114]) );
  BUF_X4 U1256 ( .A(Row2[97]), .Z(Output_1Row2[97]) );
  BUF_X4 U1257 ( .A(Row2[113]), .Z(Output_1Row2[113]) );
  BUF_X4 U1258 ( .A(Row2[9]), .Z(Output_1Row2[9]) );
  BUF_X4 U1259 ( .A(Row2[25]), .Z(Output_1Row2[25]) );
  BUF_X4 U1260 ( .A(Row2[8]), .Z(Output_1Row2[8]) );
  BUF_X4 U1261 ( .A(Row2[24]), .Z(Output_1Row2[24]) );
  BUF_X4 U1262 ( .A(Row2[7]), .Z(Output_1Row2[7]) );
  BUF_X4 U1263 ( .A(Row2[23]), .Z(Output_1Row2[23]) );
  BUF_X4 U1264 ( .A(Row2[6]), .Z(Output_1Row2[6]) );
  BUF_X4 U1265 ( .A(Row2[22]), .Z(Output_1Row2[22]) );
  BUF_X4 U1266 ( .A(Row2[5]), .Z(Output_1Row2[5]) );
  BUF_X4 U1267 ( .A(Row2[21]), .Z(Output_1Row2[21]) );
  BUF_X4 U1268 ( .A(Row2[4]), .Z(Output_1Row2[4]) );
  BUF_X4 U1269 ( .A(Row2[20]), .Z(Output_1Row2[20]) );
  BUF_X4 U1270 ( .A(Row2[3]), .Z(Output_1Row2[3]) );
  BUF_X4 U1271 ( .A(Row2[19]), .Z(Output_1Row2[19]) );
  BUF_X4 U1272 ( .A(Row2[2]), .Z(Output_1Row2[2]) );
  BUF_X4 U1273 ( .A(Row2[18]), .Z(Output_1Row2[18]) );
  BUF_X4 U1274 ( .A(Row2[1]), .Z(Output_1Row2[1]) );
  BUF_X4 U1275 ( .A(Row2[17]), .Z(Output_1Row2[17]) );
  BUF_X4 U1276 ( .A(Row1[9]), .Z(Output_1Row1[9]) );
  BUF_X4 U1277 ( .A(Row1[25]), .Z(Output_1Row1[25]) );
  BUF_X4 U1278 ( .A(Row1[8]), .Z(Output_1Row1[8]) );
  BUF_X4 U1279 ( .A(Row1[24]), .Z(Output_1Row1[24]) );
  BUF_X4 U1280 ( .A(Row1[7]), .Z(Output_1Row1[7]) );
  BUF_X4 U1281 ( .A(Row1[23]), .Z(Output_1Row1[23]) );
  BUF_X4 U1282 ( .A(Row1[6]), .Z(Output_1Row1[6]) );
  BUF_X4 U1283 ( .A(Row1[22]), .Z(Output_1Row1[22]) );
  BUF_X4 U1284 ( .A(Row1[5]), .Z(Output_1Row1[5]) );
  BUF_X4 U1285 ( .A(Row1[21]), .Z(Output_1Row1[21]) );
  BUF_X4 U1286 ( .A(Row1[4]), .Z(Output_1Row1[4]) );
  BUF_X4 U1287 ( .A(Row1[20]), .Z(Output_1Row1[20]) );
  BUF_X4 U1288 ( .A(Row1[3]), .Z(Output_1Row1[3]) );
  BUF_X4 U1289 ( .A(Row1[19]), .Z(Output_1Row1[19]) );
  BUF_X4 U1290 ( .A(Row1[2]), .Z(Output_1Row1[2]) );
  BUF_X4 U1291 ( .A(Row1[18]), .Z(Output_1Row1[18]) );
  BUF_X4 U1292 ( .A(Row1[1]), .Z(Output_1Row1[1]) );
  BUF_X4 U1293 ( .A(Row1[17]), .Z(Output_1Row1[17]) );
  BUF_X4 U1294 ( .A(Row2[169]), .Z(Output_1Row2[169]) );
  BUF_X4 U1295 ( .A(Row2[185]), .Z(Output_1Row2[185]) );
  BUF_X4 U1296 ( .A(Row2[41]), .Z(Output_1Row2[41]) );
  BUF_X4 U1297 ( .A(Row2[57]), .Z(Output_1Row2[57]) );
  BUF_X4 U1298 ( .A(Row2[168]), .Z(Output_1Row2[168]) );
  BUF_X4 U1299 ( .A(Row2[184]), .Z(Output_1Row2[184]) );
  BUF_X4 U1300 ( .A(Row2[40]), .Z(Output_1Row2[40]) );
  BUF_X4 U1301 ( .A(Row2[56]), .Z(Output_1Row2[56]) );
  BUF_X4 U1302 ( .A(Row2[167]), .Z(Output_1Row2[167]) );
  BUF_X4 U1303 ( .A(Row2[183]), .Z(Output_1Row2[183]) );
  BUF_X4 U1304 ( .A(Row2[39]), .Z(Output_1Row2[39]) );
  BUF_X4 U1305 ( .A(Row2[55]), .Z(Output_1Row2[55]) );
  BUF_X4 U1306 ( .A(Row2[166]), .Z(Output_1Row2[166]) );
  BUF_X4 U1307 ( .A(Row2[182]), .Z(Output_1Row2[182]) );
  BUF_X4 U1308 ( .A(Row2[38]), .Z(Output_1Row2[38]) );
  BUF_X4 U1309 ( .A(Row2[54]), .Z(Output_1Row2[54]) );
  BUF_X4 U1310 ( .A(Row2[165]), .Z(Output_1Row2[165]) );
  BUF_X4 U1311 ( .A(Row2[181]), .Z(Output_1Row2[181]) );
  BUF_X4 U1312 ( .A(Row2[37]), .Z(Output_1Row2[37]) );
  BUF_X4 U1313 ( .A(Row2[53]), .Z(Output_1Row2[53]) );
  BUF_X4 U1314 ( .A(Row2[164]), .Z(Output_1Row2[164]) );
  BUF_X4 U1315 ( .A(Row2[180]), .Z(Output_1Row2[180]) );
  BUF_X4 U1316 ( .A(Row2[36]), .Z(Output_1Row2[36]) );
  BUF_X4 U1317 ( .A(Row2[52]), .Z(Output_1Row2[52]) );
  BUF_X4 U1318 ( .A(Row2[163]), .Z(Output_1Row2[163]) );
  BUF_X4 U1319 ( .A(Row2[179]), .Z(Output_1Row2[179]) );
  BUF_X4 U1320 ( .A(Row2[35]), .Z(Output_1Row2[35]) );
  BUF_X4 U1321 ( .A(Row2[51]), .Z(Output_1Row2[51]) );
  BUF_X4 U1322 ( .A(Row2[162]), .Z(Output_1Row2[162]) );
  BUF_X4 U1323 ( .A(Row2[178]), .Z(Output_1Row2[178]) );
  BUF_X4 U1324 ( .A(Row2[34]), .Z(Output_1Row2[34]) );
  BUF_X4 U1325 ( .A(Row2[50]), .Z(Output_1Row2[50]) );
  BUF_X4 U1326 ( .A(Row2[161]), .Z(Output_1Row2[161]) );
  BUF_X4 U1327 ( .A(Row2[177]), .Z(Output_1Row2[177]) );
  BUF_X4 U1328 ( .A(Row2[33]), .Z(Output_1Row2[33]) );
  BUF_X4 U1329 ( .A(Row2[49]), .Z(Output_1Row2[49]) );
  BUF_X4 U1330 ( .A(Row1[169]), .Z(Output_1Row1[169]) );
  BUF_X4 U1331 ( .A(Row1[185]), .Z(Output_1Row1[185]) );
  BUF_X4 U1332 ( .A(Row1[41]), .Z(Output_1Row1[41]) );
  BUF_X4 U1333 ( .A(Row1[57]), .Z(Output_1Row1[57]) );
  BUF_X4 U1334 ( .A(Row1[168]), .Z(Output_1Row1[168]) );
  BUF_X4 U1335 ( .A(Row1[184]), .Z(Output_1Row1[184]) );
  BUF_X4 U1336 ( .A(Row1[40]), .Z(Output_1Row1[40]) );
  BUF_X4 U1337 ( .A(Row1[56]), .Z(Output_1Row1[56]) );
  BUF_X4 U1338 ( .A(Row1[167]), .Z(Output_1Row1[167]) );
  BUF_X4 U1339 ( .A(Row1[183]), .Z(Output_1Row1[183]) );
  BUF_X4 U1340 ( .A(Row1[39]), .Z(Output_1Row1[39]) );
  BUF_X4 U1341 ( .A(Row1[55]), .Z(Output_1Row1[55]) );
  BUF_X4 U1342 ( .A(Row1[166]), .Z(Output_1Row1[166]) );
  BUF_X4 U1343 ( .A(Row1[182]), .Z(Output_1Row1[182]) );
  BUF_X4 U1344 ( .A(Row1[38]), .Z(Output_1Row1[38]) );
  BUF_X4 U1345 ( .A(Row1[54]), .Z(Output_1Row1[54]) );
  BUF_X4 U1346 ( .A(Row1[165]), .Z(Output_1Row1[165]) );
  BUF_X4 U1347 ( .A(Row1[181]), .Z(Output_1Row1[181]) );
  BUF_X4 U1348 ( .A(Row1[37]), .Z(Output_1Row1[37]) );
  BUF_X4 U1349 ( .A(Row1[53]), .Z(Output_1Row1[53]) );
  BUF_X4 U1350 ( .A(Row1[164]), .Z(Output_1Row1[164]) );
  BUF_X4 U1351 ( .A(Row1[180]), .Z(Output_1Row1[180]) );
  BUF_X4 U1352 ( .A(Row1[36]), .Z(Output_1Row1[36]) );
  BUF_X4 U1353 ( .A(Row1[52]), .Z(Output_1Row1[52]) );
  BUF_X4 U1354 ( .A(Row1[163]), .Z(Output_1Row1[163]) );
  BUF_X4 U1355 ( .A(Row1[179]), .Z(Output_1Row1[179]) );
  BUF_X4 U1356 ( .A(Row1[35]), .Z(Output_1Row1[35]) );
  BUF_X4 U1357 ( .A(Row1[51]), .Z(Output_1Row1[51]) );
  BUF_X4 U1358 ( .A(Row1[162]), .Z(Output_1Row1[162]) );
  BUF_X4 U1359 ( .A(Row1[178]), .Z(Output_1Row1[178]) );
  BUF_X4 U1360 ( .A(Row1[34]), .Z(Output_1Row1[34]) );
  BUF_X4 U1361 ( .A(Row1[50]), .Z(Output_1Row1[50]) );
  BUF_X4 U1362 ( .A(Row1[161]), .Z(Output_1Row1[161]) );
  BUF_X4 U1363 ( .A(Row1[177]), .Z(Output_1Row1[177]) );
  BUF_X4 U1364 ( .A(Row1[33]), .Z(Output_1Row1[33]) );
  BUF_X4 U1365 ( .A(Row1[49]), .Z(Output_1Row1[49]) );
  BUF_X4 U1366 ( .A(PaddedRow[128]), .Z(WriteBus[128]) );
  BUF_X4 U1367 ( .A(Row1[128]), .Z(OutputPaddedRow[128]) );
  BUF_X4 U1368 ( .A(PaddedRow[129]), .Z(WriteBus[129]) );
  BUF_X4 U1369 ( .A(Row1[129]), .Z(OutputPaddedRow[129]) );
  BUF_X4 U1370 ( .A(PaddedRow[130]), .Z(WriteBus[130]) );
  BUF_X4 U1371 ( .A(Row1[130]), .Z(OutputPaddedRow[130]) );
  BUF_X4 U1372 ( .A(PaddedRow[131]), .Z(WriteBus[131]) );
  BUF_X4 U1373 ( .A(Row1[131]), .Z(OutputPaddedRow[131]) );
  BUF_X4 U1374 ( .A(PaddedRow[132]), .Z(WriteBus[132]) );
  BUF_X4 U1375 ( .A(Row1[132]), .Z(OutputPaddedRow[132]) );
  BUF_X4 U1376 ( .A(PaddedRow[133]), .Z(WriteBus[133]) );
  BUF_X4 U1377 ( .A(Row1[133]), .Z(OutputPaddedRow[133]) );
  BUF_X4 U1378 ( .A(PaddedRow[134]), .Z(WriteBus[134]) );
  BUF_X4 U1379 ( .A(Row1[134]), .Z(OutputPaddedRow[134]) );
  BUF_X4 U1380 ( .A(PaddedRow[135]), .Z(WriteBus[135]) );
  BUF_X4 U1381 ( .A(Row1[135]), .Z(OutputPaddedRow[135]) );
  BUF_X4 U1382 ( .A(PaddedRow[136]), .Z(WriteBus[136]) );
  BUF_X4 U1383 ( .A(Row1[136]), .Z(OutputPaddedRow[136]) );
  BUF_X4 U1384 ( .A(PaddedRow[137]), .Z(WriteBus[137]) );
  BUF_X4 U1385 ( .A(Row1[137]), .Z(OutputPaddedRow[137]) );
  BUF_X4 U1386 ( .A(PaddedRow[138]), .Z(WriteBus[138]) );
  BUF_X4 U1387 ( .A(Row1[138]), .Z(OutputPaddedRow[138]) );
  BUF_X4 U1388 ( .A(PaddedRow[139]), .Z(WriteBus[139]) );
  BUF_X4 U1389 ( .A(Row1[139]), .Z(OutputPaddedRow[139]) );
  BUF_X4 U1390 ( .A(PaddedRow[140]), .Z(WriteBus[140]) );
  BUF_X4 U1391 ( .A(Row1[140]), .Z(OutputPaddedRow[140]) );
  BUF_X4 U1392 ( .A(PaddedRow[141]), .Z(WriteBus[141]) );
  BUF_X4 U1393 ( .A(Row1[141]), .Z(OutputPaddedRow[141]) );
  BUF_X4 U1394 ( .A(PaddedRow[142]), .Z(WriteBus[142]) );
  BUF_X4 U1395 ( .A(Row1[142]), .Z(OutputPaddedRow[142]) );
  BUF_X4 U1396 ( .A(PaddedRow[143]), .Z(WriteBus[143]) );
  BUF_X4 U1397 ( .A(Row1[143]), .Z(OutputPaddedRow[143]) );
  BUF_X4 U1398 ( .A(PaddedRow[144]), .Z(WriteBus[144]) );
  BUF_X4 U1399 ( .A(Row1[144]), .Z(OutputPaddedRow[144]) );
  BUF_X4 U1400 ( .A(PaddedRow[145]), .Z(WriteBus[145]) );
  BUF_X4 U1401 ( .A(Row1[145]), .Z(OutputPaddedRow[145]) );
  BUF_X4 U1402 ( .A(PaddedRow[146]), .Z(WriteBus[146]) );
  BUF_X4 U1403 ( .A(Row1[146]), .Z(OutputPaddedRow[146]) );
  BUF_X4 U1404 ( .A(PaddedRow[147]), .Z(WriteBus[147]) );
  BUF_X4 U1405 ( .A(Row1[147]), .Z(OutputPaddedRow[147]) );
  BUF_X4 U1406 ( .A(PaddedRow[148]), .Z(WriteBus[148]) );
  BUF_X4 U1407 ( .A(Row1[148]), .Z(OutputPaddedRow[148]) );
  BUF_X4 U1408 ( .A(PaddedRow[149]), .Z(WriteBus[149]) );
  BUF_X4 U1409 ( .A(Row1[149]), .Z(OutputPaddedRow[149]) );
  BUF_X4 U1410 ( .A(PaddedRow[150]), .Z(WriteBus[150]) );
  BUF_X4 U1411 ( .A(Row1[150]), .Z(OutputPaddedRow[150]) );
  BUF_X4 U1412 ( .A(PaddedRow[151]), .Z(WriteBus[151]) );
  BUF_X4 U1413 ( .A(Row1[151]), .Z(OutputPaddedRow[151]) );
  BUF_X4 U1414 ( .A(PaddedRow[152]), .Z(WriteBus[152]) );
  BUF_X4 U1415 ( .A(Row1[152]), .Z(OutputPaddedRow[152]) );
  BUF_X4 U1416 ( .A(PaddedRow[153]), .Z(WriteBus[153]) );
  BUF_X4 U1417 ( .A(Row1[153]), .Z(OutputPaddedRow[153]) );
  BUF_X4 U1418 ( .A(PaddedRow[154]), .Z(WriteBus[154]) );
  BUF_X4 U1419 ( .A(Row1[154]), .Z(OutputPaddedRow[154]) );
  BUF_X4 U1420 ( .A(PaddedRow[155]), .Z(WriteBus[155]) );
  BUF_X4 U1421 ( .A(Row1[155]), .Z(OutputPaddedRow[155]) );
  BUF_X4 U1422 ( .A(PaddedRow[156]), .Z(WriteBus[156]) );
  BUF_X4 U1423 ( .A(Row1[156]), .Z(OutputPaddedRow[156]) );
  BUF_X4 U1424 ( .A(PaddedRow[157]), .Z(WriteBus[157]) );
  BUF_X4 U1425 ( .A(Row1[157]), .Z(OutputPaddedRow[157]) );
  BUF_X4 U1426 ( .A(PaddedRow[158]), .Z(WriteBus[158]) );
  BUF_X4 U1427 ( .A(Row1[158]), .Z(OutputPaddedRow[158]) );
  BUF_X4 U1428 ( .A(PaddedRow[159]), .Z(WriteBus[159]) );
  BUF_X4 U1429 ( .A(Row1[159]), .Z(OutputPaddedRow[159]) );
  BUF_X4 U1430 ( .A(PaddedRow[160]), .Z(WriteBus[160]) );
  BUF_X4 U1431 ( .A(Row1[160]), .Z(OutputPaddedRow[160]) );
  BUF_X4 U1432 ( .A(PaddedRow[161]), .Z(WriteBus[161]) );
  BUF_X4 U1433 ( .A(Row1[161]), .Z(OutputPaddedRow[161]) );
  BUF_X4 U1434 ( .A(PaddedRow[162]), .Z(WriteBus[162]) );
  BUF_X4 U1435 ( .A(Row1[162]), .Z(OutputPaddedRow[162]) );
  BUF_X4 U1436 ( .A(PaddedRow[163]), .Z(WriteBus[163]) );
  BUF_X4 U1437 ( .A(Row1[163]), .Z(OutputPaddedRow[163]) );
  BUF_X4 U1438 ( .A(PaddedRow[164]), .Z(WriteBus[164]) );
  BUF_X4 U1439 ( .A(Row1[164]), .Z(OutputPaddedRow[164]) );
  BUF_X4 U1440 ( .A(PaddedRow[165]), .Z(WriteBus[165]) );
  BUF_X4 U1441 ( .A(Row1[165]), .Z(OutputPaddedRow[165]) );
  BUF_X4 U1442 ( .A(PaddedRow[166]), .Z(WriteBus[166]) );
  BUF_X4 U1443 ( .A(Row1[166]), .Z(OutputPaddedRow[166]) );
  BUF_X4 U1444 ( .A(PaddedRow[167]), .Z(WriteBus[167]) );
  BUF_X4 U1445 ( .A(Row1[167]), .Z(OutputPaddedRow[167]) );
  BUF_X4 U1446 ( .A(PaddedRow[168]), .Z(WriteBus[168]) );
  BUF_X4 U1447 ( .A(Row1[168]), .Z(OutputPaddedRow[168]) );
  BUF_X4 U1448 ( .A(PaddedRow[169]), .Z(WriteBus[169]) );
  BUF_X4 U1449 ( .A(Row1[169]), .Z(OutputPaddedRow[169]) );
  BUF_X4 U1450 ( .A(PaddedRow[170]), .Z(WriteBus[170]) );
  BUF_X4 U1451 ( .A(Row1[170]), .Z(OutputPaddedRow[170]) );
  BUF_X4 U1452 ( .A(PaddedRow[171]), .Z(WriteBus[171]) );
  BUF_X4 U1453 ( .A(Row1[171]), .Z(OutputPaddedRow[171]) );
  BUF_X4 U1454 ( .A(PaddedRow[172]), .Z(WriteBus[172]) );
  BUF_X4 U1455 ( .A(Row1[172]), .Z(OutputPaddedRow[172]) );
  BUF_X4 U1456 ( .A(PaddedRow[173]), .Z(WriteBus[173]) );
  BUF_X4 U1457 ( .A(Row1[173]), .Z(OutputPaddedRow[173]) );
  BUF_X4 U1458 ( .A(PaddedRow[174]), .Z(WriteBus[174]) );
  BUF_X4 U1459 ( .A(Row1[174]), .Z(OutputPaddedRow[174]) );
  BUF_X4 U1460 ( .A(PaddedRow[175]), .Z(WriteBus[175]) );
  BUF_X4 U1461 ( .A(Row1[175]), .Z(OutputPaddedRow[175]) );
  BUF_X4 U1462 ( .A(Row2[111]), .Z(Output_2Row2[111]) );
  BUF_X4 U1463 ( .A(Row2[64]), .Z(Output_2Row2[64]) );
  BUF_X4 U1464 ( .A(Row2[65]), .Z(Output_2Row2[65]) );
  BUF_X4 U1465 ( .A(Row2[66]), .Z(Output_2Row2[66]) );
  BUF_X4 U1466 ( .A(Row2[67]), .Z(Output_2Row2[67]) );
  BUF_X4 U1467 ( .A(Row2[68]), .Z(Output_2Row2[68]) );
  BUF_X4 U1468 ( .A(Row2[69]), .Z(Output_2Row2[69]) );
  BUF_X4 U1469 ( .A(Row2[70]), .Z(Output_2Row2[70]) );
  BUF_X4 U1470 ( .A(Row2[71]), .Z(Output_2Row2[71]) );
  BUF_X4 U1471 ( .A(Row2[72]), .Z(Output_2Row2[72]) );
  BUF_X4 U1472 ( .A(Row2[73]), .Z(Output_2Row2[73]) );
  BUF_X4 U1473 ( .A(Row2[74]), .Z(Output_2Row2[74]) );
  BUF_X4 U1474 ( .A(Row2[75]), .Z(Output_2Row2[75]) );
  BUF_X4 U1475 ( .A(Row2[76]), .Z(Output_2Row2[76]) );
  BUF_X4 U1476 ( .A(Row2[77]), .Z(Output_2Row2[77]) );
  BUF_X4 U1477 ( .A(Row2[78]), .Z(Output_2Row2[78]) );
  BUF_X4 U1478 ( .A(Row2[79]), .Z(Output_2Row2[79]) );
  BUF_X4 U1479 ( .A(Row2[80]), .Z(Output_2Row2[80]) );
  BUF_X4 U1480 ( .A(Row2[81]), .Z(Output_2Row2[81]) );
  BUF_X4 U1481 ( .A(Row2[82]), .Z(Output_2Row2[82]) );
  BUF_X4 U1482 ( .A(Row2[83]), .Z(Output_2Row2[83]) );
  BUF_X4 U1483 ( .A(Row2[84]), .Z(Output_2Row2[84]) );
  BUF_X4 U1484 ( .A(Row2[85]), .Z(Output_2Row2[85]) );
  BUF_X4 U1485 ( .A(Row2[86]), .Z(Output_2Row2[86]) );
  BUF_X4 U1486 ( .A(Row2[87]), .Z(Output_2Row2[87]) );
  BUF_X4 U1487 ( .A(Row2[88]), .Z(Output_2Row2[88]) );
  BUF_X4 U1488 ( .A(Row2[89]), .Z(Output_2Row2[89]) );
  BUF_X4 U1489 ( .A(Row2[90]), .Z(Output_2Row2[90]) );
  BUF_X4 U1490 ( .A(Row2[91]), .Z(Output_2Row2[91]) );
  BUF_X4 U1491 ( .A(Row2[92]), .Z(Output_2Row2[92]) );
  BUF_X4 U1492 ( .A(Row2[93]), .Z(Output_2Row2[93]) );
  BUF_X4 U1493 ( .A(Row2[94]), .Z(Output_2Row2[94]) );
  BUF_X4 U1494 ( .A(Row2[95]), .Z(Output_2Row2[95]) );
  BUF_X4 U1495 ( .A(Row2[96]), .Z(Output_2Row2[96]) );
  BUF_X4 U1496 ( .A(Row2[97]), .Z(Output_2Row2[97]) );
  BUF_X4 U1497 ( .A(Row2[98]), .Z(Output_2Row2[98]) );
  BUF_X4 U1498 ( .A(Row2[99]), .Z(Output_2Row2[99]) );
  BUF_X4 U1499 ( .A(Row2[100]), .Z(Output_2Row2[100]) );
  BUF_X4 U1500 ( .A(Row2[101]), .Z(Output_2Row2[101]) );
  BUF_X4 U1501 ( .A(Row2[102]), .Z(Output_2Row2[102]) );
  BUF_X4 U1502 ( .A(Row2[103]), .Z(Output_2Row2[103]) );
  BUF_X4 U1503 ( .A(Row2[104]), .Z(Output_2Row2[104]) );
  BUF_X4 U1504 ( .A(Row2[105]), .Z(Output_2Row2[105]) );
  BUF_X4 U1505 ( .A(Row2[106]), .Z(Output_2Row2[106]) );
  BUF_X4 U1506 ( .A(Row2[107]), .Z(Output_2Row2[107]) );
  BUF_X4 U1507 ( .A(Row2[108]), .Z(Output_2Row2[108]) );
  BUF_X4 U1508 ( .A(Row2[109]), .Z(Output_2Row2[109]) );
  BUF_X4 U1509 ( .A(Row2[110]), .Z(Output_2Row2[110]) );
  BUF_X4 U1510 ( .A(Row2[47]), .Z(Output_2Row2[47]) );
  BUF_X4 U1511 ( .A(Row2[175]), .Z(Output_2Row2[175]) );
  BUF_X4 U1512 ( .A(Row2[128]), .Z(Output_2Row2[128]) );
  BUF_X4 U1513 ( .A(Row2[129]), .Z(Output_2Row2[129]) );
  BUF_X4 U1514 ( .A(Row2[130]), .Z(Output_2Row2[130]) );
  BUF_X4 U1515 ( .A(Row2[131]), .Z(Output_2Row2[131]) );
  BUF_X4 U1516 ( .A(Row2[132]), .Z(Output_2Row2[132]) );
  BUF_X4 U1517 ( .A(Row2[133]), .Z(Output_2Row2[133]) );
  BUF_X4 U1518 ( .A(Row2[134]), .Z(Output_2Row2[134]) );
  BUF_X4 U1519 ( .A(Row2[135]), .Z(Output_2Row2[135]) );
  BUF_X4 U1520 ( .A(Row2[136]), .Z(Output_2Row2[136]) );
  BUF_X4 U1521 ( .A(Row2[137]), .Z(Output_2Row2[137]) );
  BUF_X4 U1522 ( .A(Row2[138]), .Z(Output_2Row2[138]) );
  BUF_X4 U1523 ( .A(Row2[139]), .Z(Output_2Row2[139]) );
  BUF_X4 U1524 ( .A(Row2[140]), .Z(Output_2Row2[140]) );
  BUF_X4 U1525 ( .A(Row2[141]), .Z(Output_2Row2[141]) );
  BUF_X4 U1526 ( .A(Row2[142]), .Z(Output_2Row2[142]) );
  BUF_X4 U1527 ( .A(Row2[143]), .Z(Output_2Row2[143]) );
  BUF_X4 U1528 ( .A(Row2[144]), .Z(Output_2Row2[144]) );
  BUF_X4 U1529 ( .A(Row2[145]), .Z(Output_2Row2[145]) );
  BUF_X4 U1530 ( .A(Row2[146]), .Z(Output_2Row2[146]) );
  BUF_X4 U1531 ( .A(Row2[147]), .Z(Output_2Row2[147]) );
  BUF_X4 U1532 ( .A(Row2[148]), .Z(Output_2Row2[148]) );
  BUF_X4 U1533 ( .A(Row2[149]), .Z(Output_2Row2[149]) );
  BUF_X4 U1534 ( .A(Row2[150]), .Z(Output_2Row2[150]) );
  BUF_X4 U1535 ( .A(Row2[151]), .Z(Output_2Row2[151]) );
  BUF_X4 U1536 ( .A(Row2[152]), .Z(Output_2Row2[152]) );
  BUF_X4 U1537 ( .A(Row2[153]), .Z(Output_2Row2[153]) );
  BUF_X4 U1538 ( .A(Row2[154]), .Z(Output_2Row2[154]) );
  BUF_X4 U1539 ( .A(Row2[155]), .Z(Output_2Row2[155]) );
  BUF_X4 U1540 ( .A(Row2[156]), .Z(Output_2Row2[156]) );
  BUF_X4 U1541 ( .A(Row2[157]), .Z(Output_2Row2[157]) );
  BUF_X4 U1542 ( .A(Row2[158]), .Z(Output_2Row2[158]) );
  BUF_X4 U1543 ( .A(Row2[159]), .Z(Output_2Row2[159]) );
  BUF_X4 U1544 ( .A(Row2[160]), .Z(Output_2Row2[160]) );
  BUF_X4 U1545 ( .A(Row2[161]), .Z(Output_2Row2[161]) );
  BUF_X4 U1546 ( .A(Row2[162]), .Z(Output_2Row2[162]) );
  BUF_X4 U1547 ( .A(Row2[163]), .Z(Output_2Row2[163]) );
  BUF_X4 U1548 ( .A(Row2[164]), .Z(Output_2Row2[164]) );
  BUF_X4 U1549 ( .A(Row2[165]), .Z(Output_2Row2[165]) );
  BUF_X4 U1550 ( .A(Row2[166]), .Z(Output_2Row2[166]) );
  BUF_X4 U1551 ( .A(Row2[167]), .Z(Output_2Row2[167]) );
  BUF_X4 U1552 ( .A(Row2[168]), .Z(Output_2Row2[168]) );
  BUF_X4 U1553 ( .A(Row2[169]), .Z(Output_2Row2[169]) );
  BUF_X4 U1554 ( .A(Row2[170]), .Z(Output_2Row2[170]) );
  BUF_X4 U1555 ( .A(Row2[171]), .Z(Output_2Row2[171]) );
  BUF_X4 U1556 ( .A(Row2[172]), .Z(Output_2Row2[172]) );
  BUF_X4 U1557 ( .A(Row2[173]), .Z(Output_2Row2[173]) );
  BUF_X4 U1558 ( .A(Row2[174]), .Z(Output_2Row2[174]) );
  BUF_X4 U1559 ( .A(Row2[0]), .Z(Output_2Row2[0]) );
  BUF_X4 U1560 ( .A(Row2[1]), .Z(Output_2Row2[1]) );
  BUF_X4 U1561 ( .A(Row2[2]), .Z(Output_2Row2[2]) );
  BUF_X4 U1562 ( .A(Row2[3]), .Z(Output_2Row2[3]) );
  BUF_X4 U1563 ( .A(Row2[4]), .Z(Output_2Row2[4]) );
  BUF_X4 U1564 ( .A(Row2[5]), .Z(Output_2Row2[5]) );
  BUF_X4 U1565 ( .A(Row2[6]), .Z(Output_2Row2[6]) );
  BUF_X4 U1566 ( .A(Row2[7]), .Z(Output_2Row2[7]) );
  BUF_X4 U1567 ( .A(Row2[8]), .Z(Output_2Row2[8]) );
  BUF_X4 U1568 ( .A(Row2[9]), .Z(Output_2Row2[9]) );
  BUF_X4 U1569 ( .A(Row2[10]), .Z(Output_2Row2[10]) );
  BUF_X4 U1570 ( .A(Row2[11]), .Z(Output_2Row2[11]) );
  BUF_X4 U1571 ( .A(Row2[12]), .Z(Output_2Row2[12]) );
  BUF_X4 U1572 ( .A(Row2[13]), .Z(Output_2Row2[13]) );
  BUF_X4 U1573 ( .A(Row2[14]), .Z(Output_2Row2[14]) );
  BUF_X4 U1574 ( .A(Row2[15]), .Z(Output_2Row2[15]) );
  BUF_X4 U1575 ( .A(Row2[16]), .Z(Output_2Row2[16]) );
  BUF_X4 U1576 ( .A(Row2[17]), .Z(Output_2Row2[17]) );
  BUF_X4 U1577 ( .A(Row2[18]), .Z(Output_2Row2[18]) );
  BUF_X4 U1578 ( .A(Row2[19]), .Z(Output_2Row2[19]) );
  BUF_X4 U1579 ( .A(Row2[20]), .Z(Output_2Row2[20]) );
  BUF_X4 U1580 ( .A(Row2[21]), .Z(Output_2Row2[21]) );
  BUF_X4 U1581 ( .A(Row2[22]), .Z(Output_2Row2[22]) );
  BUF_X4 U1582 ( .A(Row2[23]), .Z(Output_2Row2[23]) );
  BUF_X4 U1583 ( .A(Row2[24]), .Z(Output_2Row2[24]) );
  BUF_X4 U1584 ( .A(Row2[25]), .Z(Output_2Row2[25]) );
  BUF_X4 U1585 ( .A(Row2[26]), .Z(Output_2Row2[26]) );
  BUF_X4 U1586 ( .A(Row2[27]), .Z(Output_2Row2[27]) );
  BUF_X4 U1587 ( .A(Row2[28]), .Z(Output_2Row2[28]) );
  BUF_X4 U1588 ( .A(Row2[29]), .Z(Output_2Row2[29]) );
  BUF_X4 U1589 ( .A(Row2[30]), .Z(Output_2Row2[30]) );
  BUF_X4 U1590 ( .A(Row2[31]), .Z(Output_2Row2[31]) );
  BUF_X4 U1591 ( .A(Row2[32]), .Z(Output_2Row2[32]) );
  BUF_X4 U1592 ( .A(Row2[33]), .Z(Output_2Row2[33]) );
  BUF_X4 U1593 ( .A(Row2[34]), .Z(Output_2Row2[34]) );
  BUF_X4 U1594 ( .A(Row2[35]), .Z(Output_2Row2[35]) );
  BUF_X4 U1595 ( .A(Row2[36]), .Z(Output_2Row2[36]) );
  BUF_X4 U1596 ( .A(Row2[37]), .Z(Output_2Row2[37]) );
  BUF_X4 U1597 ( .A(Row2[38]), .Z(Output_2Row2[38]) );
  BUF_X4 U1598 ( .A(Row2[39]), .Z(Output_2Row2[39]) );
  BUF_X4 U1599 ( .A(Row2[40]), .Z(Output_2Row2[40]) );
  BUF_X4 U1600 ( .A(Row2[41]), .Z(Output_2Row2[41]) );
  BUF_X4 U1601 ( .A(Row2[42]), .Z(Output_2Row2[42]) );
  BUF_X4 U1602 ( .A(Row2[43]), .Z(Output_2Row2[43]) );
  BUF_X4 U1603 ( .A(Row2[44]), .Z(Output_2Row2[44]) );
  BUF_X4 U1604 ( .A(Row2[45]), .Z(Output_2Row2[45]) );
  BUF_X4 U1605 ( .A(Row2[46]), .Z(Output_2Row2[46]) );
  BUF_X4 U1606 ( .A(Row1[192]), .Z(Output_2Row1[192]) );
  BUF_X4 U1607 ( .A(Row1[193]), .Z(Output_2Row1[193]) );
  BUF_X4 U1608 ( .A(Row1[194]), .Z(Output_2Row1[194]) );
  BUF_X4 U1609 ( .A(Row1[195]), .Z(Output_2Row1[195]) );
  BUF_X4 U1610 ( .A(Row1[196]), .Z(Output_2Row1[196]) );
  BUF_X4 U1611 ( .A(Row1[197]), .Z(Output_2Row1[197]) );
  BUF_X4 U1612 ( .A(Row1[198]), .Z(Output_2Row1[198]) );
  BUF_X4 U1613 ( .A(Row1[199]), .Z(Output_2Row1[199]) );
  BUF_X4 U1614 ( .A(Row1[200]), .Z(Output_2Row1[200]) );
  BUF_X4 U1615 ( .A(Row1[201]), .Z(Output_2Row1[201]) );
  BUF_X4 U1616 ( .A(Row1[202]), .Z(Output_2Row1[202]) );
  BUF_X4 U1617 ( .A(Row1[203]), .Z(Output_2Row1[203]) );
  BUF_X4 U1618 ( .A(Row1[204]), .Z(Output_2Row1[204]) );
  BUF_X4 U1619 ( .A(Row1[205]), .Z(Output_2Row1[205]) );
  BUF_X4 U1620 ( .A(Row1[206]), .Z(Output_2Row1[206]) );
  BUF_X4 U1621 ( .A(Row1[207]), .Z(Output_2Row1[207]) );
  BUF_X4 U1622 ( .A(Row1[208]), .Z(Output_2Row1[208]) );
  BUF_X4 U1623 ( .A(Row1[209]), .Z(Output_2Row1[209]) );
  BUF_X4 U1624 ( .A(Row1[210]), .Z(Output_2Row1[210]) );
  BUF_X4 U1625 ( .A(Row1[211]), .Z(Output_2Row1[211]) );
  BUF_X4 U1626 ( .A(Row1[212]), .Z(Output_2Row1[212]) );
  BUF_X4 U1627 ( .A(Row1[213]), .Z(Output_2Row1[213]) );
  BUF_X4 U1628 ( .A(Row1[214]), .Z(Output_2Row1[214]) );
  BUF_X4 U1629 ( .A(Row1[215]), .Z(Output_2Row1[215]) );
  BUF_X4 U1630 ( .A(Row1[216]), .Z(Output_2Row1[216]) );
  BUF_X4 U1631 ( .A(Row1[217]), .Z(Output_2Row1[217]) );
  BUF_X4 U1632 ( .A(Row1[218]), .Z(Output_2Row1[218]) );
  BUF_X4 U1633 ( .A(Row1[219]), .Z(Output_2Row1[219]) );
  BUF_X4 U1634 ( .A(Row1[220]), .Z(Output_2Row1[220]) );
  BUF_X4 U1635 ( .A(Row1[221]), .Z(Output_2Row1[221]) );
  BUF_X4 U1636 ( .A(Row1[222]), .Z(Output_2Row1[222]) );
  BUF_X4 U1637 ( .A(Row1[223]), .Z(Output_2Row1[223]) );
  BUF_X4 U1638 ( .A(Row1[224]), .Z(Output_2Row1[224]) );
  BUF_X4 U1639 ( .A(Row1[225]), .Z(Output_2Row1[225]) );
  BUF_X4 U1640 ( .A(Row1[226]), .Z(Output_2Row1[226]) );
  BUF_X4 U1641 ( .A(Row1[227]), .Z(Output_2Row1[227]) );
  BUF_X4 U1642 ( .A(Row1[228]), .Z(Output_2Row1[228]) );
  BUF_X4 U1643 ( .A(Row1[229]), .Z(Output_2Row1[229]) );
  BUF_X4 U1644 ( .A(Row1[230]), .Z(Output_2Row1[230]) );
  BUF_X4 U1645 ( .A(Row1[231]), .Z(Output_2Row1[231]) );
  BUF_X4 U1646 ( .A(Row1[232]), .Z(Output_2Row1[232]) );
  BUF_X4 U1647 ( .A(Row1[233]), .Z(Output_2Row1[233]) );
  BUF_X4 U1648 ( .A(Row1[234]), .Z(Output_2Row1[234]) );
  BUF_X4 U1649 ( .A(Row1[235]), .Z(Output_2Row1[235]) );
  BUF_X4 U1650 ( .A(Row1[236]), .Z(Output_2Row1[236]) );
  BUF_X4 U1651 ( .A(Row1[237]), .Z(Output_2Row1[237]) );
  BUF_X4 U1652 ( .A(Row1[238]), .Z(Output_2Row1[238]) );
  BUF_X4 U1653 ( .A(\U3/U2/Z_0 ), .Z(FlagX) );
  AOI222_X1 U1654 ( .A1(\U3/U5/DATA1_30 ), .A2(n2959), .B1(\U3/U5/DATA2_30 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_30 ), .C2(n2958), .ZN(n140) );
  AOI222_X1 U1655 ( .A1(\U3/U5/DATA1_31 ), .A2(n2959), .B1(\U3/U5/DATA2_31 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_31 ), .C2(n2958), .ZN(n139) );
  AOI222_X1 U1656 ( .A1(\U3/U5/DATA1_32 ), .A2(n2959), .B1(\U3/U5/DATA2_32 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_32 ), .C2(n2958), .ZN(n138) );
  AOI222_X1 U1657 ( .A1(\U3/U5/DATA1_33 ), .A2(n2959), .B1(\U3/U5/DATA2_33 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_33 ), .C2(n2958), .ZN(n137) );
  AOI222_X1 U1658 ( .A1(\U3/U5/DATA1_34 ), .A2(n2959), .B1(\U3/U5/DATA2_34 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_34 ), .C2(n2958), .ZN(n136) );
  AOI222_X1 U1659 ( .A1(\U3/U5/DATA1_35 ), .A2(n2959), .B1(\U3/U5/DATA2_35 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_35 ), .C2(n2958), .ZN(n135) );
  OAI211_X2 U1660 ( .C1(n1830), .C2(n48), .A(n49), .B(n37), .ZN(n47) );
  AOI222_X1 U1661 ( .A1(\U3/U5/DATA1_0 ), .A2(n2959), .B1(\U3/U5/DATA2_0 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_0 ), .C2(n2958), .ZN(n164) );
  AOI222_X1 U1662 ( .A1(\U3/U5/DATA1_1 ), .A2(n2959), .B1(\U3/U5/DATA2_1 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_1 ), .C2(n2958), .ZN(n163) );
  AOI222_X1 U1663 ( .A1(\U3/U5/DATA1_10 ), .A2(n2959), .B1(\U3/U5/DATA2_10 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_10 ), .C2(n2958), .ZN(n162) );
  AOI222_X1 U1664 ( .A1(\U3/U5/DATA1_11 ), .A2(n2959), .B1(\U3/U5/DATA2_11 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_11 ), .C2(n2958), .ZN(n161) );
  AOI222_X1 U1665 ( .A1(\U3/U5/DATA1_12 ), .A2(n2959), .B1(\U3/U5/DATA2_12 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_12 ), .C2(n2958), .ZN(n160) );
  AOI222_X1 U1666 ( .A1(\U3/U5/DATA1_13 ), .A2(n2959), .B1(\U3/U5/DATA2_13 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_13 ), .C2(n2958), .ZN(n159) );
  AOI222_X1 U1667 ( .A1(\U3/U5/DATA1_14 ), .A2(n2959), .B1(\U3/U5/DATA2_14 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_14 ), .C2(n2958), .ZN(n158) );
  AOI222_X1 U1668 ( .A1(\U3/U5/DATA1_15 ), .A2(n4768), .B1(\U3/U5/DATA2_15 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_15 ), .C2(n2958), .ZN(n157) );
  AOI222_X1 U1669 ( .A1(\U3/U5/DATA1_16 ), .A2(n4768), .B1(\U3/U5/DATA2_16 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_16 ), .C2(n2958), .ZN(n156) );
  AOI222_X1 U1670 ( .A1(\U3/U5/DATA1_17 ), .A2(n4768), .B1(\U3/U5/DATA2_17 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_17 ), .C2(n2958), .ZN(n155) );
  AOI222_X1 U1671 ( .A1(\U3/U5/DATA1_18 ), .A2(n4769), .B1(\U3/U5/DATA2_18 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_18 ), .C2(n2958), .ZN(n154) );
  AOI222_X1 U1672 ( .A1(\U3/U5/DATA1_19 ), .A2(n4769), .B1(\U3/U5/DATA2_19 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_19 ), .C2(n2958), .ZN(n153) );
  AOI222_X1 U1673 ( .A1(\U3/U5/DATA1_4 ), .A2(n2959), .B1(\U3/U5/DATA2_4 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_4 ), .C2(n2958), .ZN(n130) );
  AOI222_X1 U1674 ( .A1(\U3/U5/DATA1_5 ), .A2(n2959), .B1(\U3/U5/DATA2_5 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_5 ), .C2(n2958), .ZN(n121) );
  AOI222_X1 U1675 ( .A1(\U3/U5/DATA1_6 ), .A2(n2959), .B1(\U3/U5/DATA2_6 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_6 ), .C2(n2958), .ZN(n120) );
  AOI222_X1 U1676 ( .A1(\U3/U5/DATA1_7 ), .A2(n2959), .B1(\U3/U5/DATA2_7 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_7 ), .C2(n2958), .ZN(n119) );
  AOI222_X1 U1677 ( .A1(\U3/U5/DATA1_8 ), .A2(n2959), .B1(\U3/U5/DATA2_8 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_8 ), .C2(n2958), .ZN(n118) );
  AOI222_X1 U1678 ( .A1(\U3/U5/DATA1_9 ), .A2(n2959), .B1(\U3/U5/DATA2_9 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_9 ), .C2(n2958), .ZN(n116) );
  AOI222_X1 U1679 ( .A1(\U3/U5/DATA1_36 ), .A2(n2959), .B1(\U3/U5/DATA2_36 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_36 ), .C2(n2958), .ZN(n134) );
  AOI222_X1 U1680 ( .A1(\U3/U5/DATA1_37 ), .A2(n2959), .B1(\U3/U5/DATA2_37 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_37 ), .C2(n2958), .ZN(n133) );
  AOI222_X1 U1681 ( .A1(\U3/U5/DATA1_38 ), .A2(n2959), .B1(\U3/U5/DATA2_38 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_38 ), .C2(n2958), .ZN(n132) );
  AOI222_X1 U1682 ( .A1(\U3/U5/DATA1_39 ), .A2(n2959), .B1(\U3/U5/DATA2_39 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_39 ), .C2(n2958), .ZN(n131) );
  AOI222_X1 U1683 ( .A1(\U3/U5/DATA1_40 ), .A2(n2959), .B1(\U3/U5/DATA2_40 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_40 ), .C2(n2958), .ZN(n129) );
  AOI222_X1 U1684 ( .A1(\U3/U5/DATA1_41 ), .A2(n2959), .B1(\U3/U5/DATA2_41 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_41 ), .C2(n2958), .ZN(n128) );
  AOI222_X1 U1685 ( .A1(\U3/U5/DATA1_42 ), .A2(n2959), .B1(\U3/U5/DATA2_42 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_42 ), .C2(n2958), .ZN(n127) );
  AOI222_X1 U1686 ( .A1(\U3/U5/DATA1_43 ), .A2(n2959), .B1(\U3/U5/DATA2_43 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_43 ), .C2(n2958), .ZN(n126) );
  AOI222_X1 U1687 ( .A1(\U3/U5/DATA1_44 ), .A2(n2959), .B1(\U3/U5/DATA2_44 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_44 ), .C2(n2958), .ZN(n125) );
  AOI222_X1 U1688 ( .A1(\U3/U5/DATA1_45 ), .A2(n2959), .B1(\U3/U5/DATA2_45 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_45 ), .C2(n2958), .ZN(n124) );
  AOI222_X1 U1689 ( .A1(\U3/U5/DATA1_46 ), .A2(n2959), .B1(\U3/U5/DATA2_46 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_46 ), .C2(n2958), .ZN(n123) );
  AOI222_X1 U1690 ( .A1(\U3/U5/DATA1_47 ), .A2(n2959), .B1(\U3/U5/DATA2_47 ), 
        .B2(n4799), .C1(\U3/U5/DATA3_47 ), .C2(n2958), .ZN(n122) );
  NOR3_X2 U1691 ( .A1(n4770), .A2(n1830), .A3(n1828), .ZN(n82) );
  AOI22_X2 U1692 ( .A1(\U3/U7/DATA6_0 ), .A2(n4798), .B1(\U3/U7/DATA5_0 ), 
        .B2(n4802), .ZN(n72) );
  AOI22_X2 U1693 ( .A1(\U3/U7/DATA6_1 ), .A2(n4798), .B1(\U3/U7/DATA5_1 ), 
        .B2(n4802), .ZN(n71) );
  AOI22_X2 U1694 ( .A1(\U3/U7/DATA6_2 ), .A2(n4798), .B1(\U3/U7/DATA5_2 ), 
        .B2(n4802), .ZN(n70) );
  AOI22_X2 U1695 ( .A1(\U3/U7/DATA6_3 ), .A2(n4798), .B1(\U3/U7/DATA5_3 ), 
        .B2(n4802), .ZN(n69) );
  AOI22_X2 U1696 ( .A1(\U3/U7/DATA6_4 ), .A2(n4798), .B1(\U3/U7/DATA5_4 ), 
        .B2(n4802), .ZN(n68) );
  AOI22_X2 U1697 ( .A1(\U3/U7/DATA6_5 ), .A2(n4798), .B1(\U3/U7/DATA5_5 ), 
        .B2(n4802), .ZN(n67) );
  AOI22_X2 U1698 ( .A1(\U3/U7/DATA6_6 ), .A2(n4798), .B1(\U3/U7/DATA5_6 ), 
        .B2(n4802), .ZN(n66) );
  AOI22_X2 U1699 ( .A1(\U3/U7/DATA6_7 ), .A2(n4798), .B1(\U3/U7/DATA5_7 ), 
        .B2(n4802), .ZN(n65) );
  AOI22_X2 U1700 ( .A1(\U3/U7/DATA6_8 ), .A2(n4798), .B1(\U3/U7/DATA5_8 ), 
        .B2(n4802), .ZN(n75) );
  AOI22_X2 U1701 ( .A1(\U3/U7/DATA6_9 ), .A2(n4798), .B1(\U3/U7/DATA5_9 ), 
        .B2(n4802), .ZN(n74) );
  AOI22_X2 U1702 ( .A1(\U3/U7/DATA6_10 ), .A2(n4798), .B1(\U3/U7/DATA5_10 ), 
        .B2(n4802), .ZN(n73) );
  AOI211_X2 U1703 ( .C1(n4802), .C2(n45), .A(n4798), .B(n46), .ZN(n44) );
  AOI22_X2 U1704 ( .A1(n41), .A2(\U3/U4/DATA2_0 ), .B1(n4770), .B2(n42), .ZN(
        n40) );
  BUF_X4 U1705 ( .A(Row2[192]), .Z(Output_2Row2[192]) );
  BUF_X4 U1706 ( .A(Row2[193]), .Z(Output_2Row2[193]) );
  BUF_X4 U1707 ( .A(Row2[194]), .Z(Output_2Row2[194]) );
  BUF_X4 U1708 ( .A(Row2[195]), .Z(Output_2Row2[195]) );
  BUF_X4 U1709 ( .A(Row2[196]), .Z(Output_2Row2[196]) );
  BUF_X4 U1710 ( .A(Row2[197]), .Z(Output_2Row2[197]) );
  BUF_X4 U1711 ( .A(Row2[198]), .Z(Output_2Row2[198]) );
  BUF_X4 U1712 ( .A(Row2[199]), .Z(Output_2Row2[199]) );
  BUF_X4 U1713 ( .A(Row2[200]), .Z(Output_2Row2[200]) );
  BUF_X4 U1714 ( .A(Row2[201]), .Z(Output_2Row2[201]) );
  BUF_X4 U1715 ( .A(Row2[202]), .Z(Output_2Row2[202]) );
  BUF_X4 U1716 ( .A(Row2[203]), .Z(Output_2Row2[203]) );
  BUF_X4 U1717 ( .A(Row2[204]), .Z(Output_2Row2[204]) );
  BUF_X4 U1718 ( .A(Row2[205]), .Z(Output_2Row2[205]) );
  BUF_X4 U1719 ( .A(Row2[206]), .Z(Output_2Row2[206]) );
  BUF_X4 U1720 ( .A(Row2[207]), .Z(Output_2Row2[207]) );
  BUF_X4 U1721 ( .A(Row2[208]), .Z(Output_2Row2[208]) );
  BUF_X4 U1722 ( .A(Row2[209]), .Z(Output_2Row2[209]) );
  BUF_X4 U1723 ( .A(Row2[210]), .Z(Output_2Row2[210]) );
  BUF_X4 U1724 ( .A(Row2[211]), .Z(Output_2Row2[211]) );
  BUF_X4 U1725 ( .A(Row2[212]), .Z(Output_2Row2[212]) );
  BUF_X4 U1726 ( .A(Row2[213]), .Z(Output_2Row2[213]) );
  BUF_X4 U1727 ( .A(Row2[214]), .Z(Output_2Row2[214]) );
  BUF_X4 U1728 ( .A(Row2[215]), .Z(Output_2Row2[215]) );
  BUF_X4 U1729 ( .A(Row2[216]), .Z(Output_2Row2[216]) );
  BUF_X4 U1730 ( .A(Row2[217]), .Z(Output_2Row2[217]) );
  BUF_X4 U1731 ( .A(Row2[218]), .Z(Output_2Row2[218]) );
  BUF_X4 U1732 ( .A(Row2[219]), .Z(Output_2Row2[219]) );
  BUF_X4 U1733 ( .A(Row2[220]), .Z(Output_2Row2[220]) );
  BUF_X4 U1734 ( .A(Row2[221]), .Z(Output_2Row2[221]) );
  BUF_X4 U1735 ( .A(Row2[222]), .Z(Output_2Row2[222]) );
  BUF_X4 U1736 ( .A(Row2[223]), .Z(Output_2Row2[223]) );
  BUF_X4 U1737 ( .A(Row2[224]), .Z(Output_2Row2[224]) );
  BUF_X4 U1738 ( .A(Row2[225]), .Z(Output_2Row2[225]) );
  BUF_X4 U1739 ( .A(Row2[226]), .Z(Output_2Row2[226]) );
  BUF_X4 U1740 ( .A(Row2[227]), .Z(Output_2Row2[227]) );
  BUF_X4 U1741 ( .A(Row2[228]), .Z(Output_2Row2[228]) );
  BUF_X4 U1742 ( .A(Row2[229]), .Z(Output_2Row2[229]) );
  BUF_X4 U1743 ( .A(Row2[230]), .Z(Output_2Row2[230]) );
  BUF_X4 U1744 ( .A(Row2[231]), .Z(Output_2Row2[231]) );
  BUF_X4 U1745 ( .A(Row2[232]), .Z(Output_2Row2[232]) );
  BUF_X4 U1746 ( .A(Row2[233]), .Z(Output_2Row2[233]) );
  BUF_X4 U1747 ( .A(Row2[234]), .Z(Output_2Row2[234]) );
  BUF_X4 U1748 ( .A(Row2[235]), .Z(Output_2Row2[235]) );
  BUF_X4 U1749 ( .A(Row2[236]), .Z(Output_2Row2[236]) );
  BUF_X4 U1750 ( .A(Row2[237]), .Z(Output_2Row2[237]) );
  BUF_X4 U1751 ( .A(Row2[238]), .Z(Output_2Row2[238]) );
  BUF_X4 U1752 ( .A(Row2[239]), .Z(Output_2Row2[239]) );
  BUF_X4 U1753 ( .A(Row1[192]), .Z(OutputCompute[192]) );
  BUF_X4 U1754 ( .A(Row1[193]), .Z(OutputCompute[193]) );
  BUF_X4 U1755 ( .A(Row1[194]), .Z(OutputCompute[194]) );
  BUF_X4 U1756 ( .A(Row1[195]), .Z(OutputCompute[195]) );
  BUF_X4 U1757 ( .A(Row1[196]), .Z(OutputCompute[196]) );
  BUF_X4 U1758 ( .A(Row1[197]), .Z(OutputCompute[197]) );
  BUF_X4 U1759 ( .A(Row1[198]), .Z(OutputCompute[198]) );
  BUF_X4 U1760 ( .A(Row1[199]), .Z(OutputCompute[199]) );
  BUF_X4 U1761 ( .A(Row1[200]), .Z(OutputCompute[200]) );
  BUF_X4 U1762 ( .A(Row1[201]), .Z(OutputCompute[201]) );
  BUF_X4 U1763 ( .A(Row1[202]), .Z(OutputCompute[202]) );
  BUF_X4 U1764 ( .A(Row1[203]), .Z(OutputCompute[203]) );
  BUF_X4 U1765 ( .A(Row1[204]), .Z(OutputCompute[204]) );
  BUF_X4 U1766 ( .A(Row1[205]), .Z(OutputCompute[205]) );
  BUF_X4 U1767 ( .A(Row1[206]), .Z(OutputCompute[206]) );
  BUF_X4 U1768 ( .A(Row1[207]), .Z(OutputCompute[207]) );
  BUF_X4 U1769 ( .A(Row1[208]), .Z(OutputCompute[208]) );
  BUF_X4 U1770 ( .A(Row1[209]), .Z(OutputCompute[209]) );
  BUF_X4 U1771 ( .A(Row1[210]), .Z(OutputCompute[210]) );
  BUF_X4 U1772 ( .A(Row1[211]), .Z(OutputCompute[211]) );
  BUF_X4 U1773 ( .A(Row1[212]), .Z(OutputCompute[212]) );
  BUF_X4 U1774 ( .A(Row1[213]), .Z(OutputCompute[213]) );
  BUF_X4 U1775 ( .A(Row1[214]), .Z(OutputCompute[214]) );
  BUF_X4 U1776 ( .A(Row1[215]), .Z(OutputCompute[215]) );
  BUF_X4 U1777 ( .A(Row1[216]), .Z(OutputCompute[216]) );
  BUF_X4 U1778 ( .A(Row1[217]), .Z(OutputCompute[217]) );
  BUF_X4 U1779 ( .A(Row1[218]), .Z(OutputCompute[218]) );
  BUF_X4 U1780 ( .A(Row1[219]), .Z(OutputCompute[219]) );
  BUF_X4 U1781 ( .A(Row1[220]), .Z(OutputCompute[220]) );
  BUF_X4 U1782 ( .A(Row1[221]), .Z(OutputCompute[221]) );
  BUF_X4 U1783 ( .A(Row1[222]), .Z(OutputCompute[222]) );
  BUF_X4 U1784 ( .A(Row1[223]), .Z(OutputCompute[223]) );
  BUF_X4 U1785 ( .A(Row1[224]), .Z(OutputCompute[224]) );
  BUF_X4 U1786 ( .A(Row1[225]), .Z(OutputCompute[225]) );
  BUF_X4 U1787 ( .A(Row1[226]), .Z(OutputCompute[226]) );
  BUF_X4 U1788 ( .A(Row1[227]), .Z(OutputCompute[227]) );
  BUF_X4 U1789 ( .A(Row1[228]), .Z(OutputCompute[228]) );
  BUF_X4 U1790 ( .A(Row1[229]), .Z(OutputCompute[229]) );
  BUF_X4 U1791 ( .A(Row1[230]), .Z(OutputCompute[230]) );
  BUF_X4 U1792 ( .A(Row1[231]), .Z(OutputCompute[231]) );
  BUF_X4 U1793 ( .A(Row1[232]), .Z(OutputCompute[232]) );
  BUF_X4 U1794 ( .A(Row1[233]), .Z(OutputCompute[233]) );
  BUF_X4 U1795 ( .A(Row1[234]), .Z(OutputCompute[234]) );
  BUF_X4 U1796 ( .A(Row1[235]), .Z(OutputCompute[235]) );
  BUF_X4 U1797 ( .A(Row1[236]), .Z(OutputCompute[236]) );
  BUF_X4 U1798 ( .A(Row1[237]), .Z(OutputCompute[237]) );
  BUF_X4 U1799 ( .A(Row1[238]), .Z(OutputCompute[238]) );
  BUF_X4 U1800 ( .A(Row1[239]), .Z(OutputCompute[239]) );
  BUF_X4 U1801 ( .A(Row1[0]), .Z(OutputCompute[0]) );
  BUF_X4 U1802 ( .A(Row1[1]), .Z(OutputCompute[1]) );
  BUF_X4 U1803 ( .A(Row1[2]), .Z(OutputCompute[2]) );
  BUF_X4 U1804 ( .A(Row1[3]), .Z(OutputCompute[3]) );
  BUF_X4 U1805 ( .A(Row1[4]), .Z(OutputCompute[4]) );
  BUF_X4 U1806 ( .A(Row1[5]), .Z(OutputCompute[5]) );
  BUF_X4 U1807 ( .A(Row1[6]), .Z(OutputCompute[6]) );
  BUF_X4 U1808 ( .A(Row1[7]), .Z(OutputCompute[7]) );
  BUF_X4 U1809 ( .A(Row1[8]), .Z(OutputCompute[8]) );
  BUF_X4 U1810 ( .A(Row1[9]), .Z(OutputCompute[9]) );
  BUF_X4 U1811 ( .A(Row1[10]), .Z(OutputCompute[10]) );
  BUF_X4 U1812 ( .A(Row1[11]), .Z(OutputCompute[11]) );
  BUF_X4 U1813 ( .A(Row1[12]), .Z(OutputCompute[12]) );
  BUF_X4 U1814 ( .A(Row1[13]), .Z(OutputCompute[13]) );
  BUF_X4 U1815 ( .A(Row1[14]), .Z(OutputCompute[14]) );
  BUF_X4 U1816 ( .A(Row1[15]), .Z(OutputCompute[15]) );
  BUF_X4 U1817 ( .A(Row1[16]), .Z(OutputCompute[16]) );
  BUF_X4 U1818 ( .A(Row1[17]), .Z(OutputCompute[17]) );
  BUF_X4 U1819 ( .A(Row1[18]), .Z(OutputCompute[18]) );
  BUF_X4 U1820 ( .A(Row1[19]), .Z(OutputCompute[19]) );
  BUF_X4 U1821 ( .A(Row1[20]), .Z(OutputCompute[20]) );
  BUF_X4 U1822 ( .A(Row1[21]), .Z(OutputCompute[21]) );
  BUF_X4 U1823 ( .A(Row1[22]), .Z(OutputCompute[22]) );
  BUF_X4 U1824 ( .A(Row1[23]), .Z(OutputCompute[23]) );
  BUF_X4 U1825 ( .A(Row1[24]), .Z(OutputCompute[24]) );
  BUF_X4 U1826 ( .A(Row1[25]), .Z(OutputCompute[25]) );
  BUF_X4 U1827 ( .A(Row1[26]), .Z(OutputCompute[26]) );
  BUF_X4 U1828 ( .A(Row1[27]), .Z(OutputCompute[27]) );
  BUF_X4 U1829 ( .A(Row1[28]), .Z(OutputCompute[28]) );
  BUF_X4 U1830 ( .A(Row1[29]), .Z(OutputCompute[29]) );
  BUF_X4 U1831 ( .A(Row1[30]), .Z(OutputCompute[30]) );
  BUF_X4 U1832 ( .A(Row1[31]), .Z(OutputCompute[31]) );
  BUF_X4 U1833 ( .A(Row1[32]), .Z(OutputCompute[32]) );
  BUF_X4 U1834 ( .A(Row1[33]), .Z(OutputCompute[33]) );
  BUF_X4 U1835 ( .A(Row1[34]), .Z(OutputCompute[34]) );
  BUF_X4 U1836 ( .A(Row1[35]), .Z(OutputCompute[35]) );
  BUF_X4 U1837 ( .A(Row1[36]), .Z(OutputCompute[36]) );
  BUF_X4 U1838 ( .A(Row1[37]), .Z(OutputCompute[37]) );
  BUF_X4 U1839 ( .A(Row1[38]), .Z(OutputCompute[38]) );
  BUF_X4 U1840 ( .A(Row1[39]), .Z(OutputCompute[39]) );
  BUF_X4 U1841 ( .A(Row1[40]), .Z(OutputCompute[40]) );
  BUF_X4 U1842 ( .A(Row1[41]), .Z(OutputCompute[41]) );
  BUF_X4 U1843 ( .A(Row1[42]), .Z(OutputCompute[42]) );
  BUF_X4 U1844 ( .A(Row1[43]), .Z(OutputCompute[43]) );
  BUF_X4 U1845 ( .A(Row1[44]), .Z(OutputCompute[44]) );
  BUF_X4 U1846 ( .A(Row1[45]), .Z(OutputCompute[45]) );
  BUF_X4 U1847 ( .A(Row1[46]), .Z(OutputCompute[46]) );
  BUF_X4 U1848 ( .A(Row1[47]), .Z(OutputCompute[47]) );
  BUF_X4 U1849 ( .A(Row1[128]), .Z(OutputCompute[128]) );
  BUF_X4 U1850 ( .A(Row1[129]), .Z(OutputCompute[129]) );
  BUF_X4 U1851 ( .A(Row1[130]), .Z(OutputCompute[130]) );
  BUF_X4 U1852 ( .A(Row1[131]), .Z(OutputCompute[131]) );
  BUF_X4 U1853 ( .A(Row1[132]), .Z(OutputCompute[132]) );
  BUF_X4 U1854 ( .A(Row1[133]), .Z(OutputCompute[133]) );
  BUF_X4 U1855 ( .A(Row1[134]), .Z(OutputCompute[134]) );
  BUF_X4 U1856 ( .A(Row1[135]), .Z(OutputCompute[135]) );
  BUF_X4 U1857 ( .A(Row1[136]), .Z(OutputCompute[136]) );
  BUF_X4 U1858 ( .A(Row1[137]), .Z(OutputCompute[137]) );
  BUF_X4 U1859 ( .A(Row1[138]), .Z(OutputCompute[138]) );
  BUF_X4 U1860 ( .A(Row1[139]), .Z(OutputCompute[139]) );
  BUF_X4 U1861 ( .A(Row1[140]), .Z(OutputCompute[140]) );
  BUF_X4 U1862 ( .A(Row1[141]), .Z(OutputCompute[141]) );
  BUF_X4 U1863 ( .A(Row1[142]), .Z(OutputCompute[142]) );
  BUF_X4 U1864 ( .A(Row1[143]), .Z(OutputCompute[143]) );
  BUF_X4 U1865 ( .A(Row1[144]), .Z(OutputCompute[144]) );
  BUF_X4 U1866 ( .A(Row1[145]), .Z(OutputCompute[145]) );
  BUF_X4 U1867 ( .A(Row1[146]), .Z(OutputCompute[146]) );
  BUF_X4 U1868 ( .A(Row1[147]), .Z(OutputCompute[147]) );
  BUF_X4 U1869 ( .A(Row1[148]), .Z(OutputCompute[148]) );
  BUF_X4 U1870 ( .A(Row1[149]), .Z(OutputCompute[149]) );
  BUF_X4 U1871 ( .A(Row1[150]), .Z(OutputCompute[150]) );
  BUF_X4 U1872 ( .A(Row1[151]), .Z(OutputCompute[151]) );
  BUF_X4 U1873 ( .A(Row1[152]), .Z(OutputCompute[152]) );
  BUF_X4 U1874 ( .A(Row1[153]), .Z(OutputCompute[153]) );
  BUF_X4 U1875 ( .A(Row1[154]), .Z(OutputCompute[154]) );
  BUF_X4 U1876 ( .A(Row1[155]), .Z(OutputCompute[155]) );
  BUF_X4 U1877 ( .A(Row1[156]), .Z(OutputCompute[156]) );
  BUF_X4 U1878 ( .A(Row1[157]), .Z(OutputCompute[157]) );
  BUF_X4 U1879 ( .A(Row1[158]), .Z(OutputCompute[158]) );
  BUF_X4 U1880 ( .A(Row1[159]), .Z(OutputCompute[159]) );
  BUF_X4 U1881 ( .A(Row1[160]), .Z(OutputCompute[160]) );
  BUF_X4 U1882 ( .A(Row1[161]), .Z(OutputCompute[161]) );
  BUF_X4 U1883 ( .A(Row1[162]), .Z(OutputCompute[162]) );
  BUF_X4 U1884 ( .A(Row1[163]), .Z(OutputCompute[163]) );
  BUF_X4 U1885 ( .A(Row1[164]), .Z(OutputCompute[164]) );
  BUF_X4 U1886 ( .A(Row1[165]), .Z(OutputCompute[165]) );
  BUF_X4 U1887 ( .A(Row1[166]), .Z(OutputCompute[166]) );
  BUF_X4 U1888 ( .A(Row1[167]), .Z(OutputCompute[167]) );
  BUF_X4 U1889 ( .A(Row1[168]), .Z(OutputCompute[168]) );
  BUF_X4 U1890 ( .A(Row1[169]), .Z(OutputCompute[169]) );
  BUF_X4 U1891 ( .A(Row1[170]), .Z(OutputCompute[170]) );
  BUF_X4 U1892 ( .A(Row1[171]), .Z(OutputCompute[171]) );
  BUF_X4 U1893 ( .A(Row1[172]), .Z(OutputCompute[172]) );
  BUF_X4 U1894 ( .A(Row1[173]), .Z(OutputCompute[173]) );
  BUF_X4 U1895 ( .A(Row1[174]), .Z(OutputCompute[174]) );
  BUF_X4 U1896 ( .A(Row1[175]), .Z(OutputCompute[175]) );
  BUF_X4 U1897 ( .A(Row1[75]), .Z(OutputCompute[75]) );
  BUF_X4 U1898 ( .A(Row1[76]), .Z(OutputCompute[76]) );
  BUF_X4 U1899 ( .A(Row1[77]), .Z(OutputCompute[77]) );
  BUF_X4 U1900 ( .A(Row1[78]), .Z(OutputCompute[78]) );
  BUF_X4 U1901 ( .A(Row1[79]), .Z(OutputCompute[79]) );
  BUF_X4 U1902 ( .A(Row1[91]), .Z(OutputCompute[91]) );
  BUF_X4 U1903 ( .A(Row1[92]), .Z(OutputCompute[92]) );
  BUF_X4 U1904 ( .A(Row1[93]), .Z(OutputCompute[93]) );
  BUF_X4 U1905 ( .A(Row1[94]), .Z(OutputCompute[94]) );
  BUF_X4 U1906 ( .A(Row1[95]), .Z(OutputCompute[95]) );
  BUF_X4 U1907 ( .A(Row1[107]), .Z(OutputCompute[107]) );
  BUF_X4 U1908 ( .A(Row1[108]), .Z(OutputCompute[108]) );
  BUF_X4 U1909 ( .A(Row1[109]), .Z(OutputCompute[109]) );
  BUF_X4 U1910 ( .A(Row1[110]), .Z(OutputCompute[110]) );
  BUF_X4 U1911 ( .A(Row1[111]), .Z(OutputCompute[111]) );
  AOI22_X2 U1912 ( .A1(\U3/U3/DATA1_4 ), .A2(n2960), .B1(\U3/U3/DATA2_4 ), 
        .B2(n4800), .ZN(n170) );
  AOI22_X2 U1913 ( .A1(\U3/U3/DATA1_5 ), .A2(n2960), .B1(\U3/U3/DATA2_5 ), 
        .B2(n4800), .ZN(n169) );
  AOI22_X2 U1914 ( .A1(\U3/U3/DATA1_6 ), .A2(n2960), .B1(\U3/U3/DATA2_6 ), 
        .B2(n4800), .ZN(n168) );
  AOI22_X2 U1915 ( .A1(\U3/U3/DATA1_7 ), .A2(n2960), .B1(\U3/U3/DATA2_7 ), 
        .B2(n4800), .ZN(n167) );
  AOI22_X2 U1916 ( .A1(\U3/U3/DATA1_8 ), .A2(n2960), .B1(\U3/U3/DATA2_8 ), 
        .B2(n4800), .ZN(n166) );
  AOI22_X2 U1917 ( .A1(\U3/U3/DATA1_9 ), .A2(n2960), .B1(\U3/U3/DATA2_9 ), 
        .B2(n4800), .ZN(n165) );
  AOI22_X2 U1918 ( .A1(\U3/U3/DATA1_10 ), .A2(n2960), .B1(\U3/U3/DATA2_10 ), 
        .B2(n4800), .ZN(n173) );
  BUF_X4 U1919 ( .A(Row1[201]), .Z(Output_1Row1[201]) );
  BUF_X4 U1920 ( .A(Row1[233]), .Z(Output_1Row1[233]) );
  BUF_X4 U1921 ( .A(Row1[137]), .Z(Output_1Row1[137]) );
  BUF_X4 U1922 ( .A(Row1[200]), .Z(Output_1Row1[200]) );
  BUF_X4 U1923 ( .A(Row1[232]), .Z(Output_1Row1[232]) );
  BUF_X4 U1924 ( .A(Row1[136]), .Z(Output_1Row1[136]) );
  BUF_X4 U1925 ( .A(Row1[199]), .Z(Output_1Row1[199]) );
  BUF_X4 U1926 ( .A(Row1[231]), .Z(Output_1Row1[231]) );
  BUF_X4 U1927 ( .A(Row1[135]), .Z(Output_1Row1[135]) );
  BUF_X4 U1928 ( .A(Row1[198]), .Z(Output_1Row1[198]) );
  BUF_X4 U1929 ( .A(Row1[230]), .Z(Output_1Row1[230]) );
  BUF_X4 U1930 ( .A(Row1[134]), .Z(Output_1Row1[134]) );
  BUF_X4 U1931 ( .A(Row1[197]), .Z(Output_1Row1[197]) );
  BUF_X4 U1932 ( .A(Row1[229]), .Z(Output_1Row1[229]) );
  BUF_X4 U1933 ( .A(Row1[133]), .Z(Output_1Row1[133]) );
  BUF_X4 U1934 ( .A(Row1[196]), .Z(Output_1Row1[196]) );
  BUF_X4 U1935 ( .A(Row1[228]), .Z(Output_1Row1[228]) );
  BUF_X4 U1936 ( .A(Row1[132]), .Z(Output_1Row1[132]) );
  BUF_X4 U1937 ( .A(Row1[195]), .Z(Output_1Row1[195]) );
  BUF_X4 U1938 ( .A(Row1[227]), .Z(Output_1Row1[227]) );
  BUF_X4 U1939 ( .A(Row1[131]), .Z(Output_1Row1[131]) );
  BUF_X4 U1940 ( .A(Row1[194]), .Z(Output_1Row1[194]) );
  BUF_X4 U1941 ( .A(Row1[226]), .Z(Output_1Row1[226]) );
  BUF_X4 U1942 ( .A(Row1[130]), .Z(Output_1Row1[130]) );
  BUF_X4 U1943 ( .A(Row1[193]), .Z(Output_1Row1[193]) );
  BUF_X4 U1944 ( .A(Row1[225]), .Z(Output_1Row1[225]) );
  BUF_X4 U1945 ( .A(Row1[129]), .Z(Output_1Row1[129]) );
  BUF_X4 U1946 ( .A(Row1[138]), .Z(Output_1Row1[138]) );
  BUF_X4 U1947 ( .A(Row1[202]), .Z(Output_1Row1[202]) );
  BUF_X4 U1948 ( .A(Row1[234]), .Z(Output_1Row1[234]) );
  BUF_X4 U1949 ( .A(Row1[10]), .Z(Output_1Row1[10]) );
  BUF_X4 U1950 ( .A(Row2[201]), .Z(Output_1Row2[201]) );
  BUF_X4 U1951 ( .A(Row2[233]), .Z(Output_1Row2[233]) );
  BUF_X4 U1952 ( .A(Row2[137]), .Z(Output_1Row2[137]) );
  BUF_X4 U1953 ( .A(Row2[200]), .Z(Output_1Row2[200]) );
  BUF_X4 U1954 ( .A(Row2[232]), .Z(Output_1Row2[232]) );
  BUF_X4 U1955 ( .A(Row2[136]), .Z(Output_1Row2[136]) );
  BUF_X4 U1956 ( .A(Row2[199]), .Z(Output_1Row2[199]) );
  BUF_X4 U1957 ( .A(Row2[231]), .Z(Output_1Row2[231]) );
  BUF_X4 U1958 ( .A(Row2[135]), .Z(Output_1Row2[135]) );
  BUF_X4 U1959 ( .A(Row2[198]), .Z(Output_1Row2[198]) );
  BUF_X4 U1960 ( .A(Row2[230]), .Z(Output_1Row2[230]) );
  BUF_X4 U1961 ( .A(Row2[134]), .Z(Output_1Row2[134]) );
  BUF_X4 U1962 ( .A(Row2[197]), .Z(Output_1Row2[197]) );
  BUF_X4 U1963 ( .A(Row2[229]), .Z(Output_1Row2[229]) );
  BUF_X4 U1964 ( .A(Row2[133]), .Z(Output_1Row2[133]) );
  BUF_X4 U1965 ( .A(Row2[196]), .Z(Output_1Row2[196]) );
  BUF_X4 U1966 ( .A(Row2[228]), .Z(Output_1Row2[228]) );
  BUF_X4 U1967 ( .A(Row2[132]), .Z(Output_1Row2[132]) );
  BUF_X4 U1968 ( .A(Row2[195]), .Z(Output_1Row2[195]) );
  BUF_X4 U1969 ( .A(Row2[227]), .Z(Output_1Row2[227]) );
  BUF_X4 U1970 ( .A(Row2[131]), .Z(Output_1Row2[131]) );
  BUF_X4 U1971 ( .A(Row2[194]), .Z(Output_1Row2[194]) );
  BUF_X4 U1972 ( .A(Row2[226]), .Z(Output_1Row2[226]) );
  BUF_X4 U1973 ( .A(Row2[130]), .Z(Output_1Row2[130]) );
  BUF_X4 U1974 ( .A(Row2[193]), .Z(Output_1Row2[193]) );
  BUF_X4 U1975 ( .A(Row2[225]), .Z(Output_1Row2[225]) );
  BUF_X4 U1976 ( .A(Row2[129]), .Z(Output_1Row2[129]) );
  BUF_X4 U1977 ( .A(Row2[138]), .Z(Output_1Row2[138]) );
  BUF_X4 U1978 ( .A(Row2[202]), .Z(Output_1Row2[202]) );
  BUF_X4 U1979 ( .A(Row2[234]), .Z(Output_1Row2[234]) );
  BUF_X4 U1980 ( .A(Row2[10]), .Z(Output_1Row2[10]) );
  BUF_X4 U1981 ( .A(Row2[74]), .Z(Output_1Row2[74]) );
  BUF_X4 U1982 ( .A(Row2[106]), .Z(Output_1Row2[106]) );
  BUF_X4 U1983 ( .A(Row1[217]), .Z(Output_1Row1[217]) );
  BUF_X4 U1984 ( .A(Row1[153]), .Z(Output_1Row1[153]) );
  BUF_X4 U1985 ( .A(Row1[216]), .Z(Output_1Row1[216]) );
  BUF_X4 U1986 ( .A(Row1[152]), .Z(Output_1Row1[152]) );
  BUF_X4 U1987 ( .A(Row1[215]), .Z(Output_1Row1[215]) );
  BUF_X4 U1988 ( .A(Row1[151]), .Z(Output_1Row1[151]) );
  BUF_X4 U1989 ( .A(Row1[214]), .Z(Output_1Row1[214]) );
  BUF_X4 U1990 ( .A(Row1[150]), .Z(Output_1Row1[150]) );
  BUF_X4 U1991 ( .A(Row1[213]), .Z(Output_1Row1[213]) );
  BUF_X4 U1992 ( .A(Row1[149]), .Z(Output_1Row1[149]) );
  BUF_X4 U1993 ( .A(Row1[212]), .Z(Output_1Row1[212]) );
  BUF_X4 U1994 ( .A(Row1[148]), .Z(Output_1Row1[148]) );
  BUF_X4 U1995 ( .A(Row1[211]), .Z(Output_1Row1[211]) );
  BUF_X4 U1996 ( .A(Row1[147]), .Z(Output_1Row1[147]) );
  BUF_X4 U1997 ( .A(Row1[210]), .Z(Output_1Row1[210]) );
  BUF_X4 U1998 ( .A(Row1[146]), .Z(Output_1Row1[146]) );
  BUF_X4 U1999 ( .A(Row1[209]), .Z(Output_1Row1[209]) );
  BUF_X4 U2000 ( .A(Row1[145]), .Z(Output_1Row1[145]) );
  BUF_X4 U2001 ( .A(Row1[154]), .Z(Output_1Row1[154]) );
  BUF_X4 U2002 ( .A(Row1[218]), .Z(Output_1Row1[218]) );
  BUF_X4 U2003 ( .A(Row1[26]), .Z(Output_1Row1[26]) );
  BUF_X4 U2004 ( .A(Row2[217]), .Z(Output_1Row2[217]) );
  BUF_X4 U2005 ( .A(Row2[249]), .Z(Output_1Row2[249]) );
  BUF_X4 U2006 ( .A(Row2[153]), .Z(Output_1Row2[153]) );
  BUF_X4 U2007 ( .A(Row2[216]), .Z(Output_1Row2[216]) );
  BUF_X4 U2008 ( .A(Row2[248]), .Z(Output_1Row2[248]) );
  BUF_X4 U2009 ( .A(Row2[152]), .Z(Output_1Row2[152]) );
  BUF_X4 U2010 ( .A(Row2[215]), .Z(Output_1Row2[215]) );
  BUF_X4 U2011 ( .A(Row2[247]), .Z(Output_1Row2[247]) );
  BUF_X4 U2012 ( .A(Row2[151]), .Z(Output_1Row2[151]) );
  BUF_X4 U2013 ( .A(Row2[214]), .Z(Output_1Row2[214]) );
  BUF_X4 U2014 ( .A(Row2[246]), .Z(Output_1Row2[246]) );
  BUF_X4 U2015 ( .A(Row2[150]), .Z(Output_1Row2[150]) );
  BUF_X4 U2016 ( .A(Row2[213]), .Z(Output_1Row2[213]) );
  BUF_X4 U2017 ( .A(Row2[245]), .Z(Output_1Row2[245]) );
  BUF_X4 U2018 ( .A(Row2[149]), .Z(Output_1Row2[149]) );
  BUF_X4 U2019 ( .A(Row2[212]), .Z(Output_1Row2[212]) );
  BUF_X4 U2020 ( .A(Row2[244]), .Z(Output_1Row2[244]) );
  BUF_X4 U2021 ( .A(Row2[148]), .Z(Output_1Row2[148]) );
  BUF_X4 U2022 ( .A(Row2[211]), .Z(Output_1Row2[211]) );
  BUF_X4 U2023 ( .A(Row2[243]), .Z(Output_1Row2[243]) );
  BUF_X4 U2024 ( .A(Row2[147]), .Z(Output_1Row2[147]) );
  BUF_X4 U2025 ( .A(Row2[210]), .Z(Output_1Row2[210]) );
  BUF_X4 U2026 ( .A(Row2[242]), .Z(Output_1Row2[242]) );
  BUF_X4 U2027 ( .A(Row2[146]), .Z(Output_1Row2[146]) );
  BUF_X4 U2028 ( .A(Row2[209]), .Z(Output_1Row2[209]) );
  BUF_X4 U2029 ( .A(Row2[241]), .Z(Output_1Row2[241]) );
  BUF_X4 U2030 ( .A(Row2[145]), .Z(Output_1Row2[145]) );
  BUF_X4 U2031 ( .A(Row2[154]), .Z(Output_1Row2[154]) );
  BUF_X4 U2032 ( .A(Row2[218]), .Z(Output_1Row2[218]) );
  BUF_X4 U2033 ( .A(Row2[250]), .Z(Output_1Row2[250]) );
  BUF_X4 U2034 ( .A(Row2[26]), .Z(Output_1Row2[26]) );
  BUF_X4 U2035 ( .A(Row2[90]), .Z(Output_1Row2[90]) );
  BUF_X4 U2036 ( .A(Row2[122]), .Z(Output_1Row2[122]) );
  AOI22_X2 U2037 ( .A1(\U3/U3/DATA1_0 ), .A2(n2960), .B1(\U3/U3/DATA2_0 ), 
        .B2(n4800), .ZN(n175) );
  AOI22_X2 U2038 ( .A1(\U3/U3/DATA1_1 ), .A2(n2960), .B1(\U3/U3/DATA2_1 ), 
        .B2(n4800), .ZN(n174) );
  AOI22_X2 U2039 ( .A1(\U3/U3/DATA1_2 ), .A2(n2960), .B1(\U3/U3/DATA2_2 ), 
        .B2(n4800), .ZN(n172) );
  AOI22_X2 U2040 ( .A1(\U3/U3/DATA1_3 ), .A2(n2960), .B1(\U3/U3/DATA2_3 ), 
        .B2(n4800), .ZN(n171) );
  NOR2_X2 U2041 ( .A1(n4768), .A2(n8), .ZN(n83) );
  INV_X4 U2042 ( .A(n47), .ZN(n4771) );
  INV_X4 U2043 ( .A(\U3/U8/DATA4_1 ), .ZN(n4772) );
  INV_X4 U2044 ( .A(\U3/U8/DATA4_0 ), .ZN(n4773) );
  INV_X4 U2045 ( .A(\U3/U8/DATA3_1 ), .ZN(n4774) );
  INV_X4 U2046 ( .A(\U3/U8/DATA3_0 ), .ZN(n4775) );
  INV_X4 U2047 ( .A(\U3/U7/DATA3_10 ), .ZN(n4776) );
  INV_X4 U2048 ( .A(\U3/U7/DATA3_9 ), .ZN(n4777) );
  INV_X4 U2049 ( .A(\U3/U7/DATA3_8 ), .ZN(n4778) );
  INV_X4 U2050 ( .A(\U3/U7/DATA3_7 ), .ZN(n4779) );
  INV_X4 U2051 ( .A(\U3/U7/DATA3_6 ), .ZN(n4780) );
  INV_X4 U2052 ( .A(\U3/U7/DATA3_5 ), .ZN(n4781) );
  INV_X4 U2053 ( .A(\U3/U7/DATA3_4 ), .ZN(n4782) );
  INV_X4 U2054 ( .A(\U3/U7/DATA3_3 ), .ZN(n4783) );
  INV_X4 U2055 ( .A(\U3/U7/DATA3_2 ), .ZN(n4784) );
  INV_X4 U2056 ( .A(\U3/U7/DATA3_1 ), .ZN(n4785) );
  INV_X4 U2057 ( .A(\U3/U7/DATA3_0 ), .ZN(n4786) );
  INV_X4 U2058 ( .A(\U3/U7/DATA4_10 ), .ZN(n4787) );
  INV_X4 U2059 ( .A(\U3/U7/DATA4_9 ), .ZN(n4788) );
  INV_X4 U2060 ( .A(\U3/U7/DATA4_8 ), .ZN(n4789) );
  INV_X4 U2061 ( .A(\U3/U7/DATA4_7 ), .ZN(n4790) );
  INV_X4 U2062 ( .A(\U3/U7/DATA4_6 ), .ZN(n4791) );
  INV_X4 U2063 ( .A(\U3/U7/DATA4_5 ), .ZN(n4792) );
  INV_X4 U2064 ( .A(\U3/U7/DATA4_4 ), .ZN(n4793) );
  INV_X4 U2065 ( .A(\U3/U7/DATA4_3 ), .ZN(n4794) );
  INV_X4 U2066 ( .A(\U3/U7/DATA4_2 ), .ZN(n4795) );
  INV_X4 U2067 ( .A(\U3/U7/DATA4_1 ), .ZN(n4796) );
  INV_X4 U2068 ( .A(\U3/U7/DATA4_0 ), .ZN(n4797) );
  INV_X4 U2069 ( .A(n51), .ZN(n4799) );
endmodule


module update_3 ( reset, clock, X, Y, NewRowX, NewRowY, DiagonalX, DiagonalY, 
        PosDX, PosDY, DiagonalDoneX, DiagonalDoneY, Row_noX, Row_noY, 
        EnableChange );
  input [15:0] X;
  input [15:0] Y;
  input [255:0] NewRowX;
  input [255:0] NewRowY;
  output [47:0] DiagonalX;
  output [47:0] DiagonalY;
  output [12:0] PosDX;
  output [12:0] PosDY;
  input [10:0] Row_noX;
  input [10:0] Row_noY;
  input reset, clock, EnableChange;
  output DiagonalDoneX, DiagonalDoneY;
  wire   \U3/U10/DATA4_0 , \U3/U10/DATA4_1 , \U3/U10/DATA4_2 ,
         \U3/U10/DATA4_3 , \U3/U10/DATA4_4 , \U3/U10/DATA4_5 ,
         \U3/U10/DATA4_6 , \U3/U10/DATA4_7 , \U3/U10/DATA4_8 ,
         \U3/U10/DATA4_9 , \U3/U10/DATA4_10 , \U3/U10/DATA4_11 ,
         \U3/U10/DATA4_12 , \U3/U10/DATA4_13 , \U3/U10/DATA4_14 ,
         \U3/U10/DATA4_15 , \U3/U10/DATA4_16 , \U3/U10/DATA4_17 ,
         \U3/U10/DATA4_18 , \U3/U10/DATA4_19 , \U3/U10/DATA4_20 ,
         \U3/U10/DATA4_21 , \U3/U10/DATA4_22 , \U3/U10/DATA4_23 ,
         \U3/U10/DATA4_24 , \U3/U10/DATA4_25 , \U3/U10/DATA4_26 ,
         \U3/U10/DATA4_27 , \U3/U10/DATA4_28 , \U3/U10/DATA4_29 ,
         \U3/U10/DATA4_30 , \U3/U10/DATA4_31 , \U3/U10/DATA4_32 ,
         \U3/U10/DATA4_33 , \U3/U10/DATA4_34 , \U3/U10/DATA4_35 ,
         \U3/U10/DATA4_36 , \U3/U10/DATA4_37 , \U3/U10/DATA4_38 ,
         \U3/U10/DATA4_39 , \U3/U10/DATA4_40 , \U3/U10/DATA4_41 ,
         \U3/U10/DATA4_42 , \U3/U10/DATA4_43 , \U3/U10/DATA4_44 ,
         \U3/U10/DATA4_45 , \U3/U10/DATA4_46 , \U3/U10/DATA4_47 ,
         \U3/U10/DATA3_0 , \U3/U10/DATA3_1 , \U3/U10/DATA3_2 ,
         \U3/U10/DATA3_3 , \U3/U10/DATA3_4 , \U3/U10/DATA3_5 ,
         \U3/U10/DATA3_6 , \U3/U10/DATA3_7 , \U3/U10/DATA3_8 ,
         \U3/U10/DATA3_9 , \U3/U10/DATA3_10 , \U3/U10/DATA3_11 ,
         \U3/U10/DATA3_12 , \U3/U10/DATA3_13 , \U3/U10/DATA3_14 ,
         \U3/U10/DATA3_15 , \U3/U10/DATA3_16 , \U3/U10/DATA3_17 ,
         \U3/U10/DATA3_18 , \U3/U10/DATA3_19 , \U3/U10/DATA3_20 ,
         \U3/U10/DATA3_21 , \U3/U10/DATA3_22 , \U3/U10/DATA3_23 ,
         \U3/U10/DATA3_24 , \U3/U10/DATA3_25 , \U3/U10/DATA3_26 ,
         \U3/U10/DATA3_27 , \U3/U10/DATA3_28 , \U3/U10/DATA3_29 ,
         \U3/U10/DATA3_30 , \U3/U10/DATA3_31 , \U3/U10/DATA3_32 ,
         \U3/U10/DATA3_33 , \U3/U10/DATA3_34 , \U3/U10/DATA3_35 ,
         \U3/U10/DATA3_36 , \U3/U10/DATA3_37 , \U3/U10/DATA3_38 ,
         \U3/U10/DATA3_39 , \U3/U10/DATA3_40 , \U3/U10/DATA3_41 ,
         \U3/U10/DATA3_42 , \U3/U10/DATA3_43 , \U3/U10/DATA3_44 ,
         \U3/U10/DATA3_45 , \U3/U10/DATA3_46 , \U3/U10/DATA3_47 ,
         \U3/U10/DATA2_0 , \U3/U10/DATA2_1 , \U3/U10/DATA2_2 ,
         \U3/U10/DATA2_3 , \U3/U10/DATA2_4 , \U3/U10/DATA2_5 ,
         \U3/U10/DATA2_6 , \U3/U10/DATA2_7 , \U3/U10/DATA2_8 ,
         \U3/U10/DATA2_9 , \U3/U10/DATA2_10 , \U3/U10/DATA2_11 ,
         \U3/U10/DATA2_12 , \U3/U10/DATA2_13 , \U3/U10/DATA2_14 ,
         \U3/U10/DATA2_15 , \U3/U10/DATA2_16 , \U3/U10/DATA2_17 ,
         \U3/U10/DATA2_18 , \U3/U10/DATA2_19 , \U3/U10/DATA2_20 ,
         \U3/U10/DATA2_21 , \U3/U10/DATA2_22 , \U3/U10/DATA2_23 ,
         \U3/U10/DATA2_24 , \U3/U10/DATA2_25 , \U3/U10/DATA2_26 ,
         \U3/U10/DATA2_27 , \U3/U10/DATA2_28 , \U3/U10/DATA2_29 ,
         \U3/U10/DATA2_30 , \U3/U10/DATA2_31 , \U3/U10/DATA2_32 ,
         \U3/U10/DATA2_33 , \U3/U10/DATA2_34 , \U3/U10/DATA2_35 ,
         \U3/U10/DATA2_36 , \U3/U10/DATA2_37 , \U3/U10/DATA2_38 ,
         \U3/U10/DATA2_39 , \U3/U10/DATA2_40 , \U3/U10/DATA2_41 ,
         \U3/U10/DATA2_42 , \U3/U10/DATA2_43 , \U3/U10/DATA2_44 ,
         \U3/U10/DATA2_45 , \U3/U10/DATA2_46 , \U3/U10/DATA2_47 ,
         \U3/U10/DATA1_0 , \U3/U10/DATA1_1 , \U3/U10/DATA1_2 ,
         \U3/U10/DATA1_3 , \U3/U10/DATA1_4 , \U3/U10/DATA1_5 ,
         \U3/U10/DATA1_6 , \U3/U10/DATA1_7 , \U3/U10/DATA1_8 ,
         \U3/U10/DATA1_9 , \U3/U10/DATA1_10 , \U3/U10/DATA1_11 ,
         \U3/U10/DATA1_12 , \U3/U10/DATA1_13 , \U3/U10/DATA1_14 ,
         \U3/U10/DATA1_15 , \U3/U10/DATA1_16 , \U3/U10/DATA1_17 ,
         \U3/U10/DATA1_18 , \U3/U10/DATA1_19 , \U3/U10/DATA1_20 ,
         \U3/U10/DATA1_21 , \U3/U10/DATA1_22 , \U3/U10/DATA1_23 ,
         \U3/U10/DATA1_24 , \U3/U10/DATA1_25 , \U3/U10/DATA1_26 ,
         \U3/U10/DATA1_27 , \U3/U10/DATA1_28 , \U3/U10/DATA1_29 ,
         \U3/U10/DATA1_30 , \U3/U10/DATA1_31 , \U3/U10/DATA1_32 ,
         \U3/U10/DATA1_33 , \U3/U10/DATA1_34 , \U3/U10/DATA1_35 ,
         \U3/U10/DATA1_36 , \U3/U10/DATA1_37 , \U3/U10/DATA1_38 ,
         \U3/U10/DATA1_39 , \U3/U10/DATA1_40 , \U3/U10/DATA1_41 ,
         \U3/U10/DATA1_42 , \U3/U10/DATA1_43 , \U3/U10/DATA1_44 ,
         \U3/U10/DATA1_45 , \U3/U10/DATA1_46 , \U3/U10/DATA1_47 ,
         \U3/U12/DATA4_0 , \U3/U12/DATA4_1 , \U3/U12/DATA4_2 ,
         \U3/U12/DATA4_3 , \U3/U12/DATA4_4 , \U3/U12/DATA4_5 ,
         \U3/U12/DATA4_6 , \U3/U12/DATA4_7 , \U3/U12/DATA4_8 ,
         \U3/U12/DATA4_9 , \U3/U12/DATA4_10 , \U3/U12/DATA4_11 ,
         \U3/U12/DATA4_12 , \U3/U12/DATA4_13 , \U3/U12/DATA4_14 ,
         \U3/U12/DATA4_15 , \U3/U12/DATA4_16 , \U3/U12/DATA4_17 ,
         \U3/U12/DATA4_18 , \U3/U12/DATA4_19 , \U3/U12/DATA4_20 ,
         \U3/U12/DATA4_21 , \U3/U12/DATA4_22 , \U3/U12/DATA4_23 ,
         \U3/U12/DATA4_24 , \U3/U12/DATA4_25 , \U3/U12/DATA4_26 ,
         \U3/U12/DATA4_27 , \U3/U12/DATA4_28 , \U3/U12/DATA4_29 ,
         \U3/U12/DATA4_30 , \U3/U12/DATA4_31 , \U3/U12/DATA4_32 ,
         \U3/U12/DATA4_33 , \U3/U12/DATA4_34 , \U3/U12/DATA4_35 ,
         \U3/U12/DATA4_36 , \U3/U12/DATA4_37 , \U3/U12/DATA4_38 ,
         \U3/U12/DATA4_39 , \U3/U12/DATA4_40 , \U3/U12/DATA4_41 ,
         \U3/U12/DATA4_42 , \U3/U12/DATA4_43 , \U3/U12/DATA4_44 ,
         \U3/U12/DATA4_45 , \U3/U12/DATA4_46 , \U3/U12/DATA4_47 ,
         \U3/U12/DATA3_0 , \U3/U12/DATA3_1 , \U3/U12/DATA3_2 ,
         \U3/U12/DATA3_3 , \U3/U12/DATA3_4 , \U3/U12/DATA3_5 ,
         \U3/U12/DATA3_6 , \U3/U12/DATA3_7 , \U3/U12/DATA3_8 ,
         \U3/U12/DATA3_9 , \U3/U12/DATA3_10 , \U3/U12/DATA3_11 ,
         \U3/U12/DATA3_12 , \U3/U12/DATA3_13 , \U3/U12/DATA3_14 ,
         \U3/U12/DATA3_15 , \U3/U12/DATA3_16 , \U3/U12/DATA3_17 ,
         \U3/U12/DATA3_18 , \U3/U12/DATA3_19 , \U3/U12/DATA3_20 ,
         \U3/U12/DATA3_21 , \U3/U12/DATA3_22 , \U3/U12/DATA3_23 ,
         \U3/U12/DATA3_24 , \U3/U12/DATA3_25 , \U3/U12/DATA3_26 ,
         \U3/U12/DATA3_27 , \U3/U12/DATA3_28 , \U3/U12/DATA3_29 ,
         \U3/U12/DATA3_30 , \U3/U12/DATA3_31 , \U3/U12/DATA3_32 ,
         \U3/U12/DATA3_33 , \U3/U12/DATA3_34 , \U3/U12/DATA3_35 ,
         \U3/U12/DATA3_36 , \U3/U12/DATA3_37 , \U3/U12/DATA3_38 ,
         \U3/U12/DATA3_39 , \U3/U12/DATA3_40 , \U3/U12/DATA3_41 ,
         \U3/U12/DATA3_42 , \U3/U12/DATA3_43 , \U3/U12/DATA3_44 ,
         \U3/U12/DATA3_45 , \U3/U12/DATA3_46 , \U3/U12/DATA3_47 ,
         \U3/U12/DATA2_0 , \U3/U12/DATA2_1 , \U3/U12/DATA2_2 ,
         \U3/U12/DATA2_3 , \U3/U12/DATA2_4 , \U3/U12/DATA2_5 ,
         \U3/U12/DATA2_6 , \U3/U12/DATA2_7 , \U3/U12/DATA2_8 ,
         \U3/U12/DATA2_9 , \U3/U12/DATA2_10 , \U3/U12/DATA2_11 ,
         \U3/U12/DATA2_12 , \U3/U12/DATA2_13 , \U3/U12/DATA2_14 ,
         \U3/U12/DATA2_15 , \U3/U12/DATA2_16 , \U3/U12/DATA2_17 ,
         \U3/U12/DATA2_18 , \U3/U12/DATA2_19 , \U3/U12/DATA2_20 ,
         \U3/U12/DATA2_21 , \U3/U12/DATA2_22 , \U3/U12/DATA2_23 ,
         \U3/U12/DATA2_24 , \U3/U12/DATA2_25 , \U3/U12/DATA2_26 ,
         \U3/U12/DATA2_27 , \U3/U12/DATA2_28 , \U3/U12/DATA2_29 ,
         \U3/U12/DATA2_30 , \U3/U12/DATA2_31 , \U3/U12/DATA2_32 ,
         \U3/U12/DATA2_33 , \U3/U12/DATA2_34 , \U3/U12/DATA2_35 ,
         \U3/U12/DATA2_36 , \U3/U12/DATA2_37 , \U3/U12/DATA2_38 ,
         \U3/U12/DATA2_39 , \U3/U12/DATA2_40 , \U3/U12/DATA2_41 ,
         \U3/U12/DATA2_42 , \U3/U12/DATA2_43 , \U3/U12/DATA2_44 ,
         \U3/U12/DATA2_45 , \U3/U12/DATA2_46 , \U3/U12/DATA2_47 ,
         \U3/U12/DATA1_0 , \U3/U12/DATA1_1 , \U3/U12/DATA1_2 ,
         \U3/U12/DATA1_3 , \U3/U12/DATA1_4 , \U3/U12/DATA1_5 ,
         \U3/U12/DATA1_6 , \U3/U12/DATA1_7 , \U3/U12/DATA1_8 ,
         \U3/U12/DATA1_9 , \U3/U12/DATA1_10 , \U3/U12/DATA1_11 ,
         \U3/U12/DATA1_12 , \U3/U12/DATA1_13 , \U3/U12/DATA1_14 ,
         \U3/U12/DATA1_15 , \U3/U12/DATA1_16 , \U3/U12/DATA1_17 ,
         \U3/U12/DATA1_18 , \U3/U12/DATA1_19 , \U3/U12/DATA1_20 ,
         \U3/U12/DATA1_21 , \U3/U12/DATA1_22 , \U3/U12/DATA1_23 ,
         \U3/U12/DATA1_24 , \U3/U12/DATA1_25 , \U3/U12/DATA1_26 ,
         \U3/U12/DATA1_27 , \U3/U12/DATA1_28 , \U3/U12/DATA1_29 ,
         \U3/U12/DATA1_30 , \U3/U12/DATA1_31 , \U3/U12/DATA1_32 ,
         \U3/U12/DATA1_33 , \U3/U12/DATA1_34 , \U3/U12/DATA1_35 ,
         \U3/U12/DATA1_36 , \U3/U12/DATA1_37 , \U3/U12/DATA1_38 ,
         \U3/U12/DATA1_39 , \U3/U12/DATA1_40 , \U3/U12/DATA1_41 ,
         \U3/U12/DATA1_42 , \U3/U12/DATA1_43 , \U3/U12/DATA1_44 ,
         \U3/U12/DATA1_45 , \U3/U12/DATA1_46 , \U3/U12/DATA1_47 ,
         \eq_169_2/A[7] , \eq_169_2/A[6] , \eq_169_2/A[5] , \eq_169_2/A[4] ,
         \eq_169_2/A[3] , \eq_169_2/A[2] , \eq_169_2/A[1] , \eq_169_2/A[0] ,
         \eq_169_2/B[7] , \eq_169_2/B[6] , \eq_169_2/B[5] , \eq_169_2/B[4] ,
         \eq_169_2/B[3] , \eq_169_2/B[2] , \eq_169_2/B[1] , \eq_169_2/B[0] ,
         \eq_162_2/A[7] , \eq_162_2/A[6] , \eq_162_2/A[5] , \eq_162_2/A[4] ,
         \eq_162_2/A[3] , \eq_162_2/A[2] , \eq_162_2/A[1] , \eq_162_2/A[0] ,
         \eq_155_2/A[7] , \eq_155_2/A[6] , \eq_155_2/A[5] , \eq_155_2/A[4] ,
         \eq_155_2/A[3] , \eq_155_2/A[2] , \eq_155_2/A[1] , \eq_155_2/A[0] ,
         \eq_147_2/A[7] , \eq_147_2/A[6] , \eq_147_2/A[5] , \eq_147_2/A[4] ,
         \eq_147_2/A[3] , \eq_147_2/A[2] , \eq_147_2/A[1] , \eq_147_2/A[0] ,
         \eq_63_2/A[7] , \eq_63_2/A[6] , \eq_63_2/A[5] , \eq_63_2/A[4] ,
         \eq_63_2/A[3] , \eq_63_2/A[2] , \eq_63_2/A[1] , \eq_63_2/A[0] ,
         \eq_63_2/B[7] , \eq_63_2/B[6] , \eq_63_2/B[5] , \eq_63_2/B[4] ,
         \eq_63_2/B[3] , \eq_63_2/B[2] , \eq_63_2/B[1] , \eq_63_2/B[0] ,
         \eq_56_2/A[7] , \eq_56_2/A[6] , \eq_56_2/A[5] , \eq_56_2/A[4] ,
         \eq_56_2/A[3] , \eq_56_2/A[2] , \eq_56_2/A[1] , \eq_56_2/A[0] ,
         \eq_49_2/A[7] , \eq_49_2/A[6] , \eq_49_2/A[5] , \eq_49_2/A[4] ,
         \eq_49_2/A[3] , \eq_49_2/A[2] , \eq_49_2/A[1] , \eq_49_2/A[0] ,
         \eq_41_2/A[7] , \eq_41_2/A[6] , \eq_41_2/A[5] , \eq_41_2/A[4] ,
         \eq_41_2/A[3] , \eq_41_2/A[2] , \eq_41_2/A[1] , \eq_41_2/A[0] , n1,
         n13, n34, n35, n36, n37, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906;
  assign \U3/U10/DATA4_0  = NewRowX[0];
  assign \U3/U10/DATA4_1  = NewRowX[1];
  assign \U3/U10/DATA4_2  = NewRowX[2];
  assign \U3/U10/DATA4_3  = NewRowX[3];
  assign \U3/U10/DATA4_4  = NewRowX[4];
  assign \U3/U10/DATA4_5  = NewRowX[5];
  assign \U3/U10/DATA4_6  = NewRowX[6];
  assign \U3/U10/DATA4_7  = NewRowX[7];
  assign \U3/U10/DATA4_8  = NewRowX[8];
  assign \U3/U10/DATA4_9  = NewRowX[9];
  assign \U3/U10/DATA4_10  = NewRowX[10];
  assign \U3/U10/DATA4_11  = NewRowX[11];
  assign \U3/U10/DATA4_12  = NewRowX[12];
  assign \U3/U10/DATA4_13  = NewRowX[13];
  assign \U3/U10/DATA4_14  = NewRowX[14];
  assign \U3/U10/DATA4_15  = NewRowX[15];
  assign \U3/U10/DATA4_16  = NewRowX[16];
  assign \U3/U10/DATA4_17  = NewRowX[17];
  assign \U3/U10/DATA4_18  = NewRowX[18];
  assign \U3/U10/DATA4_19  = NewRowX[19];
  assign \U3/U10/DATA4_20  = NewRowX[20];
  assign \U3/U10/DATA4_21  = NewRowX[21];
  assign \U3/U10/DATA4_22  = NewRowX[22];
  assign \U3/U10/DATA4_23  = NewRowX[23];
  assign \U3/U10/DATA4_24  = NewRowX[24];
  assign \U3/U10/DATA4_25  = NewRowX[25];
  assign \U3/U10/DATA4_26  = NewRowX[26];
  assign \U3/U10/DATA4_27  = NewRowX[27];
  assign \U3/U10/DATA4_28  = NewRowX[28];
  assign \U3/U10/DATA4_29  = NewRowX[29];
  assign \U3/U10/DATA4_30  = NewRowX[30];
  assign \U3/U10/DATA4_31  = NewRowX[31];
  assign \U3/U10/DATA4_32  = NewRowX[32];
  assign \U3/U10/DATA4_33  = NewRowX[33];
  assign \U3/U10/DATA4_34  = NewRowX[34];
  assign \U3/U10/DATA4_35  = NewRowX[35];
  assign \U3/U10/DATA4_36  = NewRowX[36];
  assign \U3/U10/DATA4_37  = NewRowX[37];
  assign \U3/U10/DATA4_38  = NewRowX[38];
  assign \U3/U10/DATA4_39  = NewRowX[39];
  assign \U3/U10/DATA4_40  = NewRowX[40];
  assign \U3/U10/DATA4_41  = NewRowX[41];
  assign \U3/U10/DATA4_42  = NewRowX[42];
  assign \U3/U10/DATA4_43  = NewRowX[43];
  assign \U3/U10/DATA4_44  = NewRowX[44];
  assign \U3/U10/DATA4_45  = NewRowX[45];
  assign \U3/U10/DATA4_46  = NewRowX[46];
  assign \U3/U10/DATA4_47  = NewRowX[47];
  assign \U3/U10/DATA3_0  = NewRowX[64];
  assign \U3/U10/DATA3_1  = NewRowX[65];
  assign \U3/U10/DATA3_2  = NewRowX[66];
  assign \U3/U10/DATA3_3  = NewRowX[67];
  assign \U3/U10/DATA3_4  = NewRowX[68];
  assign \U3/U10/DATA3_5  = NewRowX[69];
  assign \U3/U10/DATA3_6  = NewRowX[70];
  assign \U3/U10/DATA3_7  = NewRowX[71];
  assign \U3/U10/DATA3_8  = NewRowX[72];
  assign \U3/U10/DATA3_9  = NewRowX[73];
  assign \U3/U10/DATA3_10  = NewRowX[74];
  assign \U3/U10/DATA3_11  = NewRowX[75];
  assign \U3/U10/DATA3_12  = NewRowX[76];
  assign \U3/U10/DATA3_13  = NewRowX[77];
  assign \U3/U10/DATA3_14  = NewRowX[78];
  assign \U3/U10/DATA3_15  = NewRowX[79];
  assign \U3/U10/DATA3_16  = NewRowX[80];
  assign \U3/U10/DATA3_17  = NewRowX[81];
  assign \U3/U10/DATA3_18  = NewRowX[82];
  assign \U3/U10/DATA3_19  = NewRowX[83];
  assign \U3/U10/DATA3_20  = NewRowX[84];
  assign \U3/U10/DATA3_21  = NewRowX[85];
  assign \U3/U10/DATA3_22  = NewRowX[86];
  assign \U3/U10/DATA3_23  = NewRowX[87];
  assign \U3/U10/DATA3_24  = NewRowX[88];
  assign \U3/U10/DATA3_25  = NewRowX[89];
  assign \U3/U10/DATA3_26  = NewRowX[90];
  assign \U3/U10/DATA3_27  = NewRowX[91];
  assign \U3/U10/DATA3_28  = NewRowX[92];
  assign \U3/U10/DATA3_29  = NewRowX[93];
  assign \U3/U10/DATA3_30  = NewRowX[94];
  assign \U3/U10/DATA3_31  = NewRowX[95];
  assign \U3/U10/DATA3_32  = NewRowX[96];
  assign \U3/U10/DATA3_33  = NewRowX[97];
  assign \U3/U10/DATA3_34  = NewRowX[98];
  assign \U3/U10/DATA3_35  = NewRowX[99];
  assign \U3/U10/DATA3_36  = NewRowX[100];
  assign \U3/U10/DATA3_37  = NewRowX[101];
  assign \U3/U10/DATA3_38  = NewRowX[102];
  assign \U3/U10/DATA3_39  = NewRowX[103];
  assign \U3/U10/DATA3_40  = NewRowX[104];
  assign \U3/U10/DATA3_41  = NewRowX[105];
  assign \U3/U10/DATA3_42  = NewRowX[106];
  assign \U3/U10/DATA3_43  = NewRowX[107];
  assign \U3/U10/DATA3_44  = NewRowX[108];
  assign \U3/U10/DATA3_45  = NewRowX[109];
  assign \U3/U10/DATA3_46  = NewRowX[110];
  assign \U3/U10/DATA3_47  = NewRowX[111];
  assign \U3/U10/DATA2_0  = NewRowX[128];
  assign \U3/U10/DATA2_1  = NewRowX[129];
  assign \U3/U10/DATA2_2  = NewRowX[130];
  assign \U3/U10/DATA2_3  = NewRowX[131];
  assign \U3/U10/DATA2_4  = NewRowX[132];
  assign \U3/U10/DATA2_5  = NewRowX[133];
  assign \U3/U10/DATA2_6  = NewRowX[134];
  assign \U3/U10/DATA2_7  = NewRowX[135];
  assign \U3/U10/DATA2_8  = NewRowX[136];
  assign \U3/U10/DATA2_9  = NewRowX[137];
  assign \U3/U10/DATA2_10  = NewRowX[138];
  assign \U3/U10/DATA2_11  = NewRowX[139];
  assign \U3/U10/DATA2_12  = NewRowX[140];
  assign \U3/U10/DATA2_13  = NewRowX[141];
  assign \U3/U10/DATA2_14  = NewRowX[142];
  assign \U3/U10/DATA2_15  = NewRowX[143];
  assign \U3/U10/DATA2_16  = NewRowX[144];
  assign \U3/U10/DATA2_17  = NewRowX[145];
  assign \U3/U10/DATA2_18  = NewRowX[146];
  assign \U3/U10/DATA2_19  = NewRowX[147];
  assign \U3/U10/DATA2_20  = NewRowX[148];
  assign \U3/U10/DATA2_21  = NewRowX[149];
  assign \U3/U10/DATA2_22  = NewRowX[150];
  assign \U3/U10/DATA2_23  = NewRowX[151];
  assign \U3/U10/DATA2_24  = NewRowX[152];
  assign \U3/U10/DATA2_25  = NewRowX[153];
  assign \U3/U10/DATA2_26  = NewRowX[154];
  assign \U3/U10/DATA2_27  = NewRowX[155];
  assign \U3/U10/DATA2_28  = NewRowX[156];
  assign \U3/U10/DATA2_29  = NewRowX[157];
  assign \U3/U10/DATA2_30  = NewRowX[158];
  assign \U3/U10/DATA2_31  = NewRowX[159];
  assign \U3/U10/DATA2_32  = NewRowX[160];
  assign \U3/U10/DATA2_33  = NewRowX[161];
  assign \U3/U10/DATA2_34  = NewRowX[162];
  assign \U3/U10/DATA2_35  = NewRowX[163];
  assign \U3/U10/DATA2_36  = NewRowX[164];
  assign \U3/U10/DATA2_37  = NewRowX[165];
  assign \U3/U10/DATA2_38  = NewRowX[166];
  assign \U3/U10/DATA2_39  = NewRowX[167];
  assign \U3/U10/DATA2_40  = NewRowX[168];
  assign \U3/U10/DATA2_41  = NewRowX[169];
  assign \U3/U10/DATA2_42  = NewRowX[170];
  assign \U3/U10/DATA2_43  = NewRowX[171];
  assign \U3/U10/DATA2_44  = NewRowX[172];
  assign \U3/U10/DATA2_45  = NewRowX[173];
  assign \U3/U10/DATA2_46  = NewRowX[174];
  assign \U3/U10/DATA2_47  = NewRowX[175];
  assign \U3/U10/DATA1_0  = NewRowX[192];
  assign \U3/U10/DATA1_1  = NewRowX[193];
  assign \U3/U10/DATA1_2  = NewRowX[194];
  assign \U3/U10/DATA1_3  = NewRowX[195];
  assign \U3/U10/DATA1_4  = NewRowX[196];
  assign \U3/U10/DATA1_5  = NewRowX[197];
  assign \U3/U10/DATA1_6  = NewRowX[198];
  assign \U3/U10/DATA1_7  = NewRowX[199];
  assign \U3/U10/DATA1_8  = NewRowX[200];
  assign \U3/U10/DATA1_9  = NewRowX[201];
  assign \U3/U10/DATA1_10  = NewRowX[202];
  assign \U3/U10/DATA1_11  = NewRowX[203];
  assign \U3/U10/DATA1_12  = NewRowX[204];
  assign \U3/U10/DATA1_13  = NewRowX[205];
  assign \U3/U10/DATA1_14  = NewRowX[206];
  assign \U3/U10/DATA1_15  = NewRowX[207];
  assign \U3/U10/DATA1_16  = NewRowX[208];
  assign \U3/U10/DATA1_17  = NewRowX[209];
  assign \U3/U10/DATA1_18  = NewRowX[210];
  assign \U3/U10/DATA1_19  = NewRowX[211];
  assign \U3/U10/DATA1_20  = NewRowX[212];
  assign \U3/U10/DATA1_21  = NewRowX[213];
  assign \U3/U10/DATA1_22  = NewRowX[214];
  assign \U3/U10/DATA1_23  = NewRowX[215];
  assign \U3/U10/DATA1_24  = NewRowX[216];
  assign \U3/U10/DATA1_25  = NewRowX[217];
  assign \U3/U10/DATA1_26  = NewRowX[218];
  assign \U3/U10/DATA1_27  = NewRowX[219];
  assign \U3/U10/DATA1_28  = NewRowX[220];
  assign \U3/U10/DATA1_29  = NewRowX[221];
  assign \U3/U10/DATA1_30  = NewRowX[222];
  assign \U3/U10/DATA1_31  = NewRowX[223];
  assign \U3/U10/DATA1_32  = NewRowX[224];
  assign \U3/U10/DATA1_33  = NewRowX[225];
  assign \U3/U10/DATA1_34  = NewRowX[226];
  assign \U3/U10/DATA1_35  = NewRowX[227];
  assign \U3/U10/DATA1_36  = NewRowX[228];
  assign \U3/U10/DATA1_37  = NewRowX[229];
  assign \U3/U10/DATA1_38  = NewRowX[230];
  assign \U3/U10/DATA1_39  = NewRowX[231];
  assign \U3/U10/DATA1_40  = NewRowX[232];
  assign \U3/U10/DATA1_41  = NewRowX[233];
  assign \U3/U10/DATA1_42  = NewRowX[234];
  assign \U3/U10/DATA1_43  = NewRowX[235];
  assign \U3/U10/DATA1_44  = NewRowX[236];
  assign \U3/U10/DATA1_45  = NewRowX[237];
  assign \U3/U10/DATA1_46  = NewRowX[238];
  assign \U3/U10/DATA1_47  = NewRowX[239];
  assign \U3/U12/DATA4_0  = NewRowY[0];
  assign \U3/U12/DATA4_1  = NewRowY[1];
  assign \U3/U12/DATA4_2  = NewRowY[2];
  assign \U3/U12/DATA4_3  = NewRowY[3];
  assign \U3/U12/DATA4_4  = NewRowY[4];
  assign \U3/U12/DATA4_5  = NewRowY[5];
  assign \U3/U12/DATA4_6  = NewRowY[6];
  assign \U3/U12/DATA4_7  = NewRowY[7];
  assign \U3/U12/DATA4_8  = NewRowY[8];
  assign \U3/U12/DATA4_9  = NewRowY[9];
  assign \U3/U12/DATA4_10  = NewRowY[10];
  assign \U3/U12/DATA4_11  = NewRowY[11];
  assign \U3/U12/DATA4_12  = NewRowY[12];
  assign \U3/U12/DATA4_13  = NewRowY[13];
  assign \U3/U12/DATA4_14  = NewRowY[14];
  assign \U3/U12/DATA4_15  = NewRowY[15];
  assign \U3/U12/DATA4_16  = NewRowY[16];
  assign \U3/U12/DATA4_17  = NewRowY[17];
  assign \U3/U12/DATA4_18  = NewRowY[18];
  assign \U3/U12/DATA4_19  = NewRowY[19];
  assign \U3/U12/DATA4_20  = NewRowY[20];
  assign \U3/U12/DATA4_21  = NewRowY[21];
  assign \U3/U12/DATA4_22  = NewRowY[22];
  assign \U3/U12/DATA4_23  = NewRowY[23];
  assign \U3/U12/DATA4_24  = NewRowY[24];
  assign \U3/U12/DATA4_25  = NewRowY[25];
  assign \U3/U12/DATA4_26  = NewRowY[26];
  assign \U3/U12/DATA4_27  = NewRowY[27];
  assign \U3/U12/DATA4_28  = NewRowY[28];
  assign \U3/U12/DATA4_29  = NewRowY[29];
  assign \U3/U12/DATA4_30  = NewRowY[30];
  assign \U3/U12/DATA4_31  = NewRowY[31];
  assign \U3/U12/DATA4_32  = NewRowY[32];
  assign \U3/U12/DATA4_33  = NewRowY[33];
  assign \U3/U12/DATA4_34  = NewRowY[34];
  assign \U3/U12/DATA4_35  = NewRowY[35];
  assign \U3/U12/DATA4_36  = NewRowY[36];
  assign \U3/U12/DATA4_37  = NewRowY[37];
  assign \U3/U12/DATA4_38  = NewRowY[38];
  assign \U3/U12/DATA4_39  = NewRowY[39];
  assign \U3/U12/DATA4_40  = NewRowY[40];
  assign \U3/U12/DATA4_41  = NewRowY[41];
  assign \U3/U12/DATA4_42  = NewRowY[42];
  assign \U3/U12/DATA4_43  = NewRowY[43];
  assign \U3/U12/DATA4_44  = NewRowY[44];
  assign \U3/U12/DATA4_45  = NewRowY[45];
  assign \U3/U12/DATA4_46  = NewRowY[46];
  assign \U3/U12/DATA4_47  = NewRowY[47];
  assign \U3/U12/DATA3_0  = NewRowY[64];
  assign \U3/U12/DATA3_1  = NewRowY[65];
  assign \U3/U12/DATA3_2  = NewRowY[66];
  assign \U3/U12/DATA3_3  = NewRowY[67];
  assign \U3/U12/DATA3_4  = NewRowY[68];
  assign \U3/U12/DATA3_5  = NewRowY[69];
  assign \U3/U12/DATA3_6  = NewRowY[70];
  assign \U3/U12/DATA3_7  = NewRowY[71];
  assign \U3/U12/DATA3_8  = NewRowY[72];
  assign \U3/U12/DATA3_9  = NewRowY[73];
  assign \U3/U12/DATA3_10  = NewRowY[74];
  assign \U3/U12/DATA3_11  = NewRowY[75];
  assign \U3/U12/DATA3_12  = NewRowY[76];
  assign \U3/U12/DATA3_13  = NewRowY[77];
  assign \U3/U12/DATA3_14  = NewRowY[78];
  assign \U3/U12/DATA3_15  = NewRowY[79];
  assign \U3/U12/DATA3_16  = NewRowY[80];
  assign \U3/U12/DATA3_17  = NewRowY[81];
  assign \U3/U12/DATA3_18  = NewRowY[82];
  assign \U3/U12/DATA3_19  = NewRowY[83];
  assign \U3/U12/DATA3_20  = NewRowY[84];
  assign \U3/U12/DATA3_21  = NewRowY[85];
  assign \U3/U12/DATA3_22  = NewRowY[86];
  assign \U3/U12/DATA3_23  = NewRowY[87];
  assign \U3/U12/DATA3_24  = NewRowY[88];
  assign \U3/U12/DATA3_25  = NewRowY[89];
  assign \U3/U12/DATA3_26  = NewRowY[90];
  assign \U3/U12/DATA3_27  = NewRowY[91];
  assign \U3/U12/DATA3_28  = NewRowY[92];
  assign \U3/U12/DATA3_29  = NewRowY[93];
  assign \U3/U12/DATA3_30  = NewRowY[94];
  assign \U3/U12/DATA3_31  = NewRowY[95];
  assign \U3/U12/DATA3_32  = NewRowY[96];
  assign \U3/U12/DATA3_33  = NewRowY[97];
  assign \U3/U12/DATA3_34  = NewRowY[98];
  assign \U3/U12/DATA3_35  = NewRowY[99];
  assign \U3/U12/DATA3_36  = NewRowY[100];
  assign \U3/U12/DATA3_37  = NewRowY[101];
  assign \U3/U12/DATA3_38  = NewRowY[102];
  assign \U3/U12/DATA3_39  = NewRowY[103];
  assign \U3/U12/DATA3_40  = NewRowY[104];
  assign \U3/U12/DATA3_41  = NewRowY[105];
  assign \U3/U12/DATA3_42  = NewRowY[106];
  assign \U3/U12/DATA3_43  = NewRowY[107];
  assign \U3/U12/DATA3_44  = NewRowY[108];
  assign \U3/U12/DATA3_45  = NewRowY[109];
  assign \U3/U12/DATA3_46  = NewRowY[110];
  assign \U3/U12/DATA3_47  = NewRowY[111];
  assign \U3/U12/DATA2_0  = NewRowY[128];
  assign \U3/U12/DATA2_1  = NewRowY[129];
  assign \U3/U12/DATA2_2  = NewRowY[130];
  assign \U3/U12/DATA2_3  = NewRowY[131];
  assign \U3/U12/DATA2_4  = NewRowY[132];
  assign \U3/U12/DATA2_5  = NewRowY[133];
  assign \U3/U12/DATA2_6  = NewRowY[134];
  assign \U3/U12/DATA2_7  = NewRowY[135];
  assign \U3/U12/DATA2_8  = NewRowY[136];
  assign \U3/U12/DATA2_9  = NewRowY[137];
  assign \U3/U12/DATA2_10  = NewRowY[138];
  assign \U3/U12/DATA2_11  = NewRowY[139];
  assign \U3/U12/DATA2_12  = NewRowY[140];
  assign \U3/U12/DATA2_13  = NewRowY[141];
  assign \U3/U12/DATA2_14  = NewRowY[142];
  assign \U3/U12/DATA2_15  = NewRowY[143];
  assign \U3/U12/DATA2_16  = NewRowY[144];
  assign \U3/U12/DATA2_17  = NewRowY[145];
  assign \U3/U12/DATA2_18  = NewRowY[146];
  assign \U3/U12/DATA2_19  = NewRowY[147];
  assign \U3/U12/DATA2_20  = NewRowY[148];
  assign \U3/U12/DATA2_21  = NewRowY[149];
  assign \U3/U12/DATA2_22  = NewRowY[150];
  assign \U3/U12/DATA2_23  = NewRowY[151];
  assign \U3/U12/DATA2_24  = NewRowY[152];
  assign \U3/U12/DATA2_25  = NewRowY[153];
  assign \U3/U12/DATA2_26  = NewRowY[154];
  assign \U3/U12/DATA2_27  = NewRowY[155];
  assign \U3/U12/DATA2_28  = NewRowY[156];
  assign \U3/U12/DATA2_29  = NewRowY[157];
  assign \U3/U12/DATA2_30  = NewRowY[158];
  assign \U3/U12/DATA2_31  = NewRowY[159];
  assign \U3/U12/DATA2_32  = NewRowY[160];
  assign \U3/U12/DATA2_33  = NewRowY[161];
  assign \U3/U12/DATA2_34  = NewRowY[162];
  assign \U3/U12/DATA2_35  = NewRowY[163];
  assign \U3/U12/DATA2_36  = NewRowY[164];
  assign \U3/U12/DATA2_37  = NewRowY[165];
  assign \U3/U12/DATA2_38  = NewRowY[166];
  assign \U3/U12/DATA2_39  = NewRowY[167];
  assign \U3/U12/DATA2_40  = NewRowY[168];
  assign \U3/U12/DATA2_41  = NewRowY[169];
  assign \U3/U12/DATA2_42  = NewRowY[170];
  assign \U3/U12/DATA2_43  = NewRowY[171];
  assign \U3/U12/DATA2_44  = NewRowY[172];
  assign \U3/U12/DATA2_45  = NewRowY[173];
  assign \U3/U12/DATA2_46  = NewRowY[174];
  assign \U3/U12/DATA2_47  = NewRowY[175];
  assign \U3/U12/DATA1_0  = NewRowY[192];
  assign \U3/U12/DATA1_1  = NewRowY[193];
  assign \U3/U12/DATA1_2  = NewRowY[194];
  assign \U3/U12/DATA1_3  = NewRowY[195];
  assign \U3/U12/DATA1_4  = NewRowY[196];
  assign \U3/U12/DATA1_5  = NewRowY[197];
  assign \U3/U12/DATA1_6  = NewRowY[198];
  assign \U3/U12/DATA1_7  = NewRowY[199];
  assign \U3/U12/DATA1_8  = NewRowY[200];
  assign \U3/U12/DATA1_9  = NewRowY[201];
  assign \U3/U12/DATA1_10  = NewRowY[202];
  assign \U3/U12/DATA1_11  = NewRowY[203];
  assign \U3/U12/DATA1_12  = NewRowY[204];
  assign \U3/U12/DATA1_13  = NewRowY[205];
  assign \U3/U12/DATA1_14  = NewRowY[206];
  assign \U3/U12/DATA1_15  = NewRowY[207];
  assign \U3/U12/DATA1_16  = NewRowY[208];
  assign \U3/U12/DATA1_17  = NewRowY[209];
  assign \U3/U12/DATA1_18  = NewRowY[210];
  assign \U3/U12/DATA1_19  = NewRowY[211];
  assign \U3/U12/DATA1_20  = NewRowY[212];
  assign \U3/U12/DATA1_21  = NewRowY[213];
  assign \U3/U12/DATA1_22  = NewRowY[214];
  assign \U3/U12/DATA1_23  = NewRowY[215];
  assign \U3/U12/DATA1_24  = NewRowY[216];
  assign \U3/U12/DATA1_25  = NewRowY[217];
  assign \U3/U12/DATA1_26  = NewRowY[218];
  assign \U3/U12/DATA1_27  = NewRowY[219];
  assign \U3/U12/DATA1_28  = NewRowY[220];
  assign \U3/U12/DATA1_29  = NewRowY[221];
  assign \U3/U12/DATA1_30  = NewRowY[222];
  assign \U3/U12/DATA1_31  = NewRowY[223];
  assign \U3/U12/DATA1_32  = NewRowY[224];
  assign \U3/U12/DATA1_33  = NewRowY[225];
  assign \U3/U12/DATA1_34  = NewRowY[226];
  assign \U3/U12/DATA1_35  = NewRowY[227];
  assign \U3/U12/DATA1_36  = NewRowY[228];
  assign \U3/U12/DATA1_37  = NewRowY[229];
  assign \U3/U12/DATA1_38  = NewRowY[230];
  assign \U3/U12/DATA1_39  = NewRowY[231];
  assign \U3/U12/DATA1_40  = NewRowY[232];
  assign \U3/U12/DATA1_41  = NewRowY[233];
  assign \U3/U12/DATA1_42  = NewRowY[234];
  assign \U3/U12/DATA1_43  = NewRowY[235];
  assign \U3/U12/DATA1_44  = NewRowY[236];
  assign \U3/U12/DATA1_45  = NewRowY[237];
  assign \U3/U12/DATA1_46  = NewRowY[238];
  assign \U3/U12/DATA1_47  = NewRowY[239];
  assign \eq_169_2/A[7]  = NewRowY[55];
  assign \eq_169_2/A[6]  = NewRowY[54];
  assign \eq_169_2/A[5]  = NewRowY[53];
  assign \eq_169_2/A[4]  = NewRowY[52];
  assign \eq_169_2/A[3]  = NewRowY[51];
  assign \eq_169_2/A[2]  = NewRowY[50];
  assign \eq_169_2/A[1]  = NewRowY[49];
  assign \eq_169_2/A[0]  = NewRowY[48];
  assign \eq_169_2/B[7]  = Y[7];
  assign \eq_169_2/B[6]  = Y[6];
  assign \eq_169_2/B[5]  = Y[5];
  assign \eq_169_2/B[4]  = Y[4];
  assign \eq_169_2/B[3]  = Y[3];
  assign \eq_169_2/B[2]  = Y[2];
  assign \eq_169_2/B[1]  = Y[1];
  assign \eq_169_2/B[0]  = Y[0];
  assign \eq_162_2/A[7]  = NewRowY[119];
  assign \eq_162_2/A[6]  = NewRowY[118];
  assign \eq_162_2/A[5]  = NewRowY[117];
  assign \eq_162_2/A[4]  = NewRowY[116];
  assign \eq_162_2/A[3]  = NewRowY[115];
  assign \eq_162_2/A[2]  = NewRowY[114];
  assign \eq_162_2/A[1]  = NewRowY[113];
  assign \eq_162_2/A[0]  = NewRowY[112];
  assign \eq_155_2/A[7]  = NewRowY[183];
  assign \eq_155_2/A[6]  = NewRowY[182];
  assign \eq_155_2/A[5]  = NewRowY[181];
  assign \eq_155_2/A[4]  = NewRowY[180];
  assign \eq_155_2/A[3]  = NewRowY[179];
  assign \eq_155_2/A[2]  = NewRowY[178];
  assign \eq_155_2/A[1]  = NewRowY[177];
  assign \eq_155_2/A[0]  = NewRowY[176];
  assign \eq_147_2/A[7]  = NewRowY[247];
  assign \eq_147_2/A[6]  = NewRowY[246];
  assign \eq_147_2/A[5]  = NewRowY[245];
  assign \eq_147_2/A[4]  = NewRowY[244];
  assign \eq_147_2/A[3]  = NewRowY[243];
  assign \eq_147_2/A[2]  = NewRowY[242];
  assign \eq_147_2/A[1]  = NewRowY[241];
  assign \eq_147_2/A[0]  = NewRowY[240];
  assign \eq_63_2/A[7]  = NewRowX[55];
  assign \eq_63_2/A[6]  = NewRowX[54];
  assign \eq_63_2/A[5]  = NewRowX[53];
  assign \eq_63_2/A[4]  = NewRowX[52];
  assign \eq_63_2/A[3]  = NewRowX[51];
  assign \eq_63_2/A[2]  = NewRowX[50];
  assign \eq_63_2/A[1]  = NewRowX[49];
  assign \eq_63_2/A[0]  = NewRowX[48];
  assign \eq_63_2/B[7]  = X[7];
  assign \eq_63_2/B[6]  = X[6];
  assign \eq_63_2/B[5]  = X[5];
  assign \eq_63_2/B[4]  = X[4];
  assign \eq_63_2/B[3]  = X[3];
  assign \eq_63_2/B[2]  = X[2];
  assign \eq_63_2/B[1]  = X[1];
  assign \eq_63_2/B[0]  = X[0];
  assign \eq_56_2/A[7]  = NewRowX[119];
  assign \eq_56_2/A[6]  = NewRowX[118];
  assign \eq_56_2/A[5]  = NewRowX[117];
  assign \eq_56_2/A[4]  = NewRowX[116];
  assign \eq_56_2/A[3]  = NewRowX[115];
  assign \eq_56_2/A[2]  = NewRowX[114];
  assign \eq_56_2/A[1]  = NewRowX[113];
  assign \eq_56_2/A[0]  = NewRowX[112];
  assign \eq_49_2/A[7]  = NewRowX[183];
  assign \eq_49_2/A[6]  = NewRowX[182];
  assign \eq_49_2/A[5]  = NewRowX[181];
  assign \eq_49_2/A[4]  = NewRowX[180];
  assign \eq_49_2/A[3]  = NewRowX[179];
  assign \eq_49_2/A[2]  = NewRowX[178];
  assign \eq_49_2/A[1]  = NewRowX[177];
  assign \eq_49_2/A[0]  = NewRowX[176];
  assign \eq_41_2/A[7]  = NewRowX[247];
  assign \eq_41_2/A[6]  = NewRowX[246];
  assign \eq_41_2/A[5]  = NewRowX[245];
  assign \eq_41_2/A[4]  = NewRowX[244];
  assign \eq_41_2/A[3]  = NewRowX[243];
  assign \eq_41_2/A[2]  = NewRowX[242];
  assign \eq_41_2/A[1]  = NewRowX[241];
  assign \eq_41_2/A[0]  = NewRowX[240];

  DFF_X1 \DiagonalX_reg[47]  ( .D(n466), .CK(clock), .Q(DiagonalX[47]) );
  DFF_X1 \DiagonalX_reg[46]  ( .D(n465), .CK(clock), .Q(DiagonalX[46]) );
  DFF_X1 \DiagonalX_reg[45]  ( .D(n464), .CK(clock), .Q(DiagonalX[45]) );
  DFF_X1 \DiagonalX_reg[44]  ( .D(n463), .CK(clock), .Q(DiagonalX[44]) );
  DFF_X1 \DiagonalX_reg[43]  ( .D(n462), .CK(clock), .Q(DiagonalX[43]) );
  DFF_X1 \DiagonalX_reg[42]  ( .D(n461), .CK(clock), .Q(DiagonalX[42]) );
  DFF_X1 \DiagonalX_reg[41]  ( .D(n460), .CK(clock), .Q(DiagonalX[41]) );
  DFF_X1 \DiagonalX_reg[40]  ( .D(n459), .CK(clock), .Q(DiagonalX[40]) );
  DFF_X1 \DiagonalX_reg[39]  ( .D(n458), .CK(clock), .Q(DiagonalX[39]) );
  DFF_X1 \DiagonalX_reg[38]  ( .D(n457), .CK(clock), .Q(DiagonalX[38]) );
  DFF_X1 \DiagonalX_reg[37]  ( .D(n456), .CK(clock), .Q(DiagonalX[37]) );
  DFF_X1 \DiagonalX_reg[36]  ( .D(n455), .CK(clock), .Q(DiagonalX[36]) );
  DFF_X1 \DiagonalX_reg[35]  ( .D(n454), .CK(clock), .Q(DiagonalX[35]) );
  DFF_X1 \DiagonalX_reg[34]  ( .D(n453), .CK(clock), .Q(DiagonalX[34]) );
  DFF_X1 \DiagonalX_reg[33]  ( .D(n452), .CK(clock), .Q(DiagonalX[33]) );
  DFF_X1 \DiagonalX_reg[32]  ( .D(n451), .CK(clock), .Q(DiagonalX[32]) );
  DFF_X1 \DiagonalX_reg[31]  ( .D(n450), .CK(clock), .Q(DiagonalX[31]) );
  DFF_X1 \DiagonalX_reg[30]  ( .D(n449), .CK(clock), .Q(DiagonalX[30]) );
  DFF_X1 \DiagonalX_reg[29]  ( .D(n448), .CK(clock), .Q(DiagonalX[29]) );
  DFF_X1 \DiagonalX_reg[28]  ( .D(n447), .CK(clock), .Q(DiagonalX[28]) );
  DFF_X1 \DiagonalX_reg[27]  ( .D(n446), .CK(clock), .Q(DiagonalX[27]) );
  DFF_X1 \DiagonalX_reg[26]  ( .D(n445), .CK(clock), .Q(DiagonalX[26]) );
  DFF_X1 \DiagonalX_reg[25]  ( .D(n444), .CK(clock), .Q(DiagonalX[25]) );
  DFF_X1 \DiagonalX_reg[24]  ( .D(n443), .CK(clock), .Q(DiagonalX[24]) );
  DFF_X1 \DiagonalX_reg[23]  ( .D(n442), .CK(clock), .Q(DiagonalX[23]) );
  DFF_X1 \DiagonalX_reg[22]  ( .D(n441), .CK(clock), .Q(DiagonalX[22]) );
  DFF_X1 \DiagonalX_reg[21]  ( .D(n440), .CK(clock), .Q(DiagonalX[21]) );
  DFF_X1 \DiagonalX_reg[20]  ( .D(n439), .CK(clock), .Q(DiagonalX[20]) );
  DFF_X1 \DiagonalX_reg[19]  ( .D(n438), .CK(clock), .Q(DiagonalX[19]) );
  DFF_X1 \DiagonalX_reg[18]  ( .D(n437), .CK(clock), .Q(DiagonalX[18]) );
  DFF_X1 \DiagonalX_reg[17]  ( .D(n436), .CK(clock), .Q(DiagonalX[17]) );
  DFF_X1 \DiagonalX_reg[16]  ( .D(n435), .CK(clock), .Q(DiagonalX[16]) );
  DFF_X1 \DiagonalX_reg[15]  ( .D(n434), .CK(clock), .Q(DiagonalX[15]) );
  DFF_X1 \DiagonalX_reg[14]  ( .D(n433), .CK(clock), .Q(DiagonalX[14]) );
  DFF_X1 \DiagonalX_reg[13]  ( .D(n432), .CK(clock), .Q(DiagonalX[13]) );
  DFF_X1 \DiagonalX_reg[12]  ( .D(n431), .CK(clock), .Q(DiagonalX[12]) );
  DFF_X1 \DiagonalX_reg[11]  ( .D(n430), .CK(clock), .Q(DiagonalX[11]) );
  DFF_X1 \DiagonalX_reg[10]  ( .D(n429), .CK(clock), .Q(DiagonalX[10]) );
  DFF_X1 \DiagonalX_reg[9]  ( .D(n428), .CK(clock), .Q(DiagonalX[9]) );
  DFF_X1 \DiagonalX_reg[8]  ( .D(n427), .CK(clock), .Q(DiagonalX[8]) );
  DFF_X1 \DiagonalX_reg[7]  ( .D(n426), .CK(clock), .Q(DiagonalX[7]) );
  DFF_X1 \DiagonalX_reg[6]  ( .D(n425), .CK(clock), .Q(DiagonalX[6]) );
  DFF_X1 \DiagonalX_reg[5]  ( .D(n424), .CK(clock), .Q(DiagonalX[5]) );
  DFF_X1 \DiagonalX_reg[4]  ( .D(n423), .CK(clock), .Q(DiagonalX[4]) );
  DFF_X1 \DiagonalX_reg[3]  ( .D(n422), .CK(clock), .Q(DiagonalX[3]) );
  DFF_X1 \DiagonalX_reg[2]  ( .D(n421), .CK(clock), .Q(DiagonalX[2]) );
  DFF_X1 \DiagonalX_reg[1]  ( .D(n420), .CK(clock), .Q(DiagonalX[1]) );
  DFF_X1 \DiagonalX_reg[0]  ( .D(n419), .CK(clock), .Q(DiagonalX[0]) );
  DFF_X1 \PosDX_reg[12]  ( .D(n877), .CK(clock), .Q(PosDX[12]) );
  DFF_X1 \PosDX_reg[11]  ( .D(n878), .CK(clock), .Q(PosDX[11]) );
  DFF_X1 \PosDX_reg[10]  ( .D(n879), .CK(clock), .Q(PosDX[10]) );
  DFF_X1 \PosDX_reg[9]  ( .D(n880), .CK(clock), .Q(PosDX[9]) );
  DFF_X1 \PosDX_reg[8]  ( .D(n881), .CK(clock), .Q(PosDX[8]) );
  DFF_X1 \PosDX_reg[7]  ( .D(n882), .CK(clock), .Q(PosDX[7]) );
  DFF_X1 \PosDX_reg[6]  ( .D(n883), .CK(clock), .Q(PosDX[6]) );
  DFF_X1 \PosDX_reg[5]  ( .D(n884), .CK(clock), .Q(PosDX[5]) );
  DFF_X1 \PosDX_reg[4]  ( .D(n885), .CK(clock), .Q(PosDX[4]) );
  DFF_X1 \PosDX_reg[3]  ( .D(n886), .CK(clock), .Q(PosDX[3]) );
  DFF_X1 \PosDX_reg[2]  ( .D(n887), .CK(clock), .Q(PosDX[2]) );
  DFF_X1 \PosDX_reg[1]  ( .D(n417), .CK(clock), .Q(PosDX[1]) );
  DFF_X1 \PosDX_reg[0]  ( .D(n416), .CK(clock), .Q(PosDX[0]) );
  DFF_X1 \DiagonalY_reg[47]  ( .D(n415), .CK(clock), .Q(DiagonalY[47]) );
  DFF_X1 \DiagonalY_reg[46]  ( .D(n414), .CK(clock), .Q(DiagonalY[46]) );
  DFF_X1 \DiagonalY_reg[45]  ( .D(n413), .CK(clock), .Q(DiagonalY[45]) );
  DFF_X1 \DiagonalY_reg[44]  ( .D(n412), .CK(clock), .Q(DiagonalY[44]) );
  DFF_X1 \DiagonalY_reg[43]  ( .D(n411), .CK(clock), .Q(DiagonalY[43]) );
  DFF_X1 \DiagonalY_reg[42]  ( .D(n410), .CK(clock), .Q(DiagonalY[42]) );
  DFF_X1 \DiagonalY_reg[41]  ( .D(n409), .CK(clock), .Q(DiagonalY[41]) );
  DFF_X1 \DiagonalY_reg[40]  ( .D(n408), .CK(clock), .Q(DiagonalY[40]) );
  DFF_X1 \DiagonalY_reg[39]  ( .D(n407), .CK(clock), .Q(DiagonalY[39]) );
  DFF_X1 \DiagonalY_reg[38]  ( .D(n406), .CK(clock), .Q(DiagonalY[38]) );
  DFF_X1 \DiagonalY_reg[37]  ( .D(n405), .CK(clock), .Q(DiagonalY[37]) );
  DFF_X1 \DiagonalY_reg[36]  ( .D(n404), .CK(clock), .Q(DiagonalY[36]) );
  DFF_X1 \DiagonalY_reg[35]  ( .D(n403), .CK(clock), .Q(DiagonalY[35]) );
  DFF_X1 \DiagonalY_reg[34]  ( .D(n402), .CK(clock), .Q(DiagonalY[34]) );
  DFF_X1 \DiagonalY_reg[33]  ( .D(n401), .CK(clock), .Q(DiagonalY[33]) );
  DFF_X1 \DiagonalY_reg[32]  ( .D(n400), .CK(clock), .Q(DiagonalY[32]) );
  DFF_X1 \DiagonalY_reg[31]  ( .D(n399), .CK(clock), .Q(DiagonalY[31]) );
  DFF_X1 \DiagonalY_reg[30]  ( .D(n398), .CK(clock), .Q(DiagonalY[30]) );
  DFF_X1 \DiagonalY_reg[29]  ( .D(n397), .CK(clock), .Q(DiagonalY[29]) );
  DFF_X1 \DiagonalY_reg[28]  ( .D(n396), .CK(clock), .Q(DiagonalY[28]) );
  DFF_X1 \DiagonalY_reg[27]  ( .D(n395), .CK(clock), .Q(DiagonalY[27]) );
  DFF_X1 \DiagonalY_reg[26]  ( .D(n394), .CK(clock), .Q(DiagonalY[26]) );
  DFF_X1 \DiagonalY_reg[25]  ( .D(n393), .CK(clock), .Q(DiagonalY[25]) );
  DFF_X1 \DiagonalY_reg[24]  ( .D(n392), .CK(clock), .Q(DiagonalY[24]) );
  DFF_X1 \DiagonalY_reg[23]  ( .D(n391), .CK(clock), .Q(DiagonalY[23]) );
  DFF_X1 \DiagonalY_reg[22]  ( .D(n390), .CK(clock), .Q(DiagonalY[22]) );
  DFF_X1 \DiagonalY_reg[21]  ( .D(n389), .CK(clock), .Q(DiagonalY[21]) );
  DFF_X1 \DiagonalY_reg[20]  ( .D(n388), .CK(clock), .Q(DiagonalY[20]) );
  DFF_X1 \DiagonalY_reg[19]  ( .D(n387), .CK(clock), .Q(DiagonalY[19]) );
  DFF_X1 \DiagonalY_reg[18]  ( .D(n386), .CK(clock), .Q(DiagonalY[18]) );
  DFF_X1 \DiagonalY_reg[17]  ( .D(n385), .CK(clock), .Q(DiagonalY[17]) );
  DFF_X1 \DiagonalY_reg[16]  ( .D(n384), .CK(clock), .Q(DiagonalY[16]) );
  DFF_X1 \DiagonalY_reg[15]  ( .D(n383), .CK(clock), .Q(DiagonalY[15]) );
  DFF_X1 \DiagonalY_reg[14]  ( .D(n382), .CK(clock), .Q(DiagonalY[14]) );
  DFF_X1 \DiagonalY_reg[13]  ( .D(n381), .CK(clock), .Q(DiagonalY[13]) );
  DFF_X1 \DiagonalY_reg[12]  ( .D(n380), .CK(clock), .Q(DiagonalY[12]) );
  DFF_X1 \DiagonalY_reg[11]  ( .D(n379), .CK(clock), .Q(DiagonalY[11]) );
  DFF_X1 \DiagonalY_reg[10]  ( .D(n378), .CK(clock), .Q(DiagonalY[10]) );
  DFF_X1 \DiagonalY_reg[9]  ( .D(n377), .CK(clock), .Q(DiagonalY[9]) );
  DFF_X1 \DiagonalY_reg[8]  ( .D(n376), .CK(clock), .Q(DiagonalY[8]) );
  DFF_X1 \DiagonalY_reg[7]  ( .D(n375), .CK(clock), .Q(DiagonalY[7]) );
  DFF_X1 \DiagonalY_reg[6]  ( .D(n374), .CK(clock), .Q(DiagonalY[6]) );
  DFF_X1 \DiagonalY_reg[5]  ( .D(n373), .CK(clock), .Q(DiagonalY[5]) );
  DFF_X1 \DiagonalY_reg[4]  ( .D(n372), .CK(clock), .Q(DiagonalY[4]) );
  DFF_X1 \DiagonalY_reg[3]  ( .D(n371), .CK(clock), .Q(DiagonalY[3]) );
  DFF_X1 \DiagonalY_reg[2]  ( .D(n370), .CK(clock), .Q(DiagonalY[2]) );
  DFF_X1 \DiagonalY_reg[1]  ( .D(n369), .CK(clock), .Q(DiagonalY[1]) );
  DFF_X1 \DiagonalY_reg[0]  ( .D(n368), .CK(clock), .Q(DiagonalY[0]) );
  DFF_X1 \PosDY_reg[12]  ( .D(n888), .CK(clock), .Q(PosDY[12]) );
  DFF_X1 \PosDY_reg[11]  ( .D(n889), .CK(clock), .Q(PosDY[11]) );
  DFF_X1 \PosDY_reg[10]  ( .D(n890), .CK(clock), .Q(PosDY[10]) );
  DFF_X1 \PosDY_reg[9]  ( .D(n891), .CK(clock), .Q(PosDY[9]) );
  DFF_X1 \PosDY_reg[8]  ( .D(n892), .CK(clock), .Q(PosDY[8]) );
  DFF_X1 \PosDY_reg[7]  ( .D(n893), .CK(clock), .Q(PosDY[7]) );
  DFF_X1 \PosDY_reg[6]  ( .D(n894), .CK(clock), .Q(PosDY[6]) );
  DFF_X1 \PosDY_reg[5]  ( .D(n895), .CK(clock), .Q(PosDY[5]) );
  DFF_X1 \PosDY_reg[4]  ( .D(n896), .CK(clock), .Q(PosDY[4]) );
  DFF_X1 \PosDY_reg[3]  ( .D(n897), .CK(clock), .Q(PosDY[3]) );
  DFF_X1 \PosDY_reg[2]  ( .D(n898), .CK(clock), .Q(PosDY[2]) );
  DFF_X1 \PosDY_reg[1]  ( .D(n366), .CK(clock), .Q(PosDY[1]) );
  DFF_X1 \PosDY_reg[0]  ( .D(n365), .CK(clock), .Q(PosDY[0]) );
  NAND2_X2 U4 ( .A1(PosDY[0]), .A2(n899), .ZN(n35) );
  NAND2_X2 U7 ( .A1(PosDY[1]), .A2(n899), .ZN(n40) );
  OAI22_X2 U20 ( .A1(n903), .A2(n901), .B1(n54), .B2(n13), .ZN(n367) );
  NAND2_X2 U21 ( .A1(n55), .A2(n56), .ZN(n368) );
  NAND2_X2 U24 ( .A1(n59), .A2(n60), .ZN(n369) );
  NAND2_X2 U27 ( .A1(n61), .A2(n62), .ZN(n370) );
  NAND2_X2 U30 ( .A1(n63), .A2(n64), .ZN(n371) );
  NAND2_X2 U33 ( .A1(n65), .A2(n66), .ZN(n372) );
  NAND2_X2 U36 ( .A1(n67), .A2(n68), .ZN(n373) );
  NAND2_X2 U39 ( .A1(n69), .A2(n70), .ZN(n374) );
  NAND2_X2 U42 ( .A1(n71), .A2(n72), .ZN(n375) );
  NAND2_X2 U45 ( .A1(n73), .A2(n74), .ZN(n376) );
  NAND2_X2 U48 ( .A1(n75), .A2(n76), .ZN(n377) );
  NAND2_X2 U51 ( .A1(n77), .A2(n78), .ZN(n378) );
  NAND2_X2 U54 ( .A1(n79), .A2(n80), .ZN(n379) );
  NAND2_X2 U57 ( .A1(n81), .A2(n82), .ZN(n380) );
  NAND2_X2 U60 ( .A1(n83), .A2(n84), .ZN(n381) );
  NAND2_X2 U63 ( .A1(n85), .A2(n86), .ZN(n382) );
  NAND2_X2 U66 ( .A1(n87), .A2(n88), .ZN(n383) );
  NAND2_X2 U69 ( .A1(n89), .A2(n90), .ZN(n384) );
  NAND2_X2 U72 ( .A1(n91), .A2(n92), .ZN(n385) );
  NAND2_X2 U75 ( .A1(n93), .A2(n94), .ZN(n386) );
  NAND2_X2 U78 ( .A1(n95), .A2(n96), .ZN(n387) );
  NAND2_X2 U81 ( .A1(n97), .A2(n98), .ZN(n388) );
  NAND2_X2 U84 ( .A1(n99), .A2(n100), .ZN(n389) );
  NAND2_X2 U87 ( .A1(n101), .A2(n102), .ZN(n390) );
  NAND2_X2 U90 ( .A1(n103), .A2(n104), .ZN(n391) );
  NAND2_X2 U93 ( .A1(n105), .A2(n106), .ZN(n392) );
  NAND2_X2 U96 ( .A1(n107), .A2(n108), .ZN(n393) );
  NAND2_X2 U99 ( .A1(n109), .A2(n110), .ZN(n394) );
  NAND2_X2 U102 ( .A1(n111), .A2(n112), .ZN(n395) );
  NAND2_X2 U105 ( .A1(n113), .A2(n114), .ZN(n396) );
  NAND2_X2 U108 ( .A1(n115), .A2(n116), .ZN(n397) );
  NAND2_X2 U111 ( .A1(n117), .A2(n118), .ZN(n398) );
  NAND2_X2 U114 ( .A1(n119), .A2(n120), .ZN(n399) );
  NAND2_X2 U117 ( .A1(n121), .A2(n122), .ZN(n400) );
  NAND2_X2 U120 ( .A1(n123), .A2(n124), .ZN(n401) );
  NAND2_X2 U123 ( .A1(n125), .A2(n126), .ZN(n402) );
  NAND2_X2 U126 ( .A1(n127), .A2(n128), .ZN(n403) );
  NAND2_X2 U129 ( .A1(n129), .A2(n130), .ZN(n404) );
  NAND2_X2 U132 ( .A1(n131), .A2(n132), .ZN(n405) );
  NAND2_X2 U135 ( .A1(n133), .A2(n134), .ZN(n406) );
  NAND2_X2 U138 ( .A1(n135), .A2(n136), .ZN(n407) );
  NAND2_X2 U141 ( .A1(n137), .A2(n138), .ZN(n408) );
  NAND2_X2 U144 ( .A1(n139), .A2(n140), .ZN(n409) );
  NAND2_X2 U147 ( .A1(n141), .A2(n142), .ZN(n410) );
  NAND2_X2 U150 ( .A1(n143), .A2(n144), .ZN(n411) );
  NAND2_X2 U153 ( .A1(n145), .A2(n146), .ZN(n412) );
  NAND2_X2 U156 ( .A1(n147), .A2(n148), .ZN(n413) );
  NAND2_X2 U159 ( .A1(n149), .A2(n150), .ZN(n414) );
  NAND2_X2 U162 ( .A1(n151), .A2(n152), .ZN(n415) );
  NAND2_X2 U168 ( .A1(n53), .A2(n154), .ZN(n54) );
  NOR3_X2 U169 ( .A1(n155), .A2(n906), .A3(n39), .ZN(n53) );
  NAND2_X2 U170 ( .A1(n153), .A2(n37), .ZN(n39) );
  NAND4_X2 U171 ( .A1(n156), .A2(n157), .A3(n158), .A4(n159), .ZN(n153) );
  NOR4_X2 U172 ( .A1(n160), .A2(n161), .A3(n162), .A4(n163), .ZN(n159) );
  XOR2_X2 U173 ( .A(\eq_169_2/B[0] ), .B(\eq_155_2/A[0] ), .Z(n163) );
  XOR2_X2 U174 ( .A(\eq_169_2/B[2] ), .B(\eq_155_2/A[2] ), .Z(n162) );
  XOR2_X2 U175 ( .A(\eq_169_2/B[1] ), .B(\eq_155_2/A[1] ), .Z(n161) );
  NAND3_X2 U176 ( .A1(NewRowY[190]), .A2(NewRowY[189]), .A3(NewRowY[191]), 
        .ZN(n160) );
  NOR3_X2 U177 ( .A1(n164), .A2(n165), .A3(n166), .ZN(n158) );
  XOR2_X2 U178 ( .A(\eq_169_2/B[3] ), .B(\eq_155_2/A[3] ), .Z(n166) );
  XOR2_X2 U179 ( .A(\eq_169_2/B[5] ), .B(\eq_155_2/A[5] ), .Z(n165) );
  XOR2_X2 U180 ( .A(\eq_169_2/B[4] ), .B(\eq_155_2/A[4] ), .Z(n164) );
  XNOR2_X2 U181 ( .A(\eq_169_2/B[6] ), .B(\eq_155_2/A[6] ), .ZN(n157) );
  XNOR2_X2 U182 ( .A(\eq_169_2/B[7] ), .B(\eq_155_2/A[7] ), .ZN(n156) );
  NAND4_X2 U183 ( .A1(n167), .A2(n168), .A3(n169), .A4(n170), .ZN(n36) );
  NOR4_X2 U184 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(n170) );
  XOR2_X2 U185 ( .A(\eq_169_2/B[0] ), .B(\eq_162_2/A[0] ), .Z(n174) );
  XOR2_X2 U186 ( .A(\eq_169_2/B[2] ), .B(\eq_162_2/A[2] ), .Z(n173) );
  XOR2_X2 U187 ( .A(\eq_169_2/B[1] ), .B(\eq_162_2/A[1] ), .Z(n172) );
  NAND3_X2 U188 ( .A1(NewRowY[126]), .A2(NewRowY[125]), .A3(NewRowY[127]), 
        .ZN(n171) );
  NOR3_X2 U189 ( .A1(n175), .A2(n176), .A3(n177), .ZN(n169) );
  XOR2_X2 U190 ( .A(\eq_169_2/B[3] ), .B(\eq_162_2/A[3] ), .Z(n177) );
  XOR2_X2 U191 ( .A(\eq_169_2/B[5] ), .B(\eq_162_2/A[5] ), .Z(n176) );
  XOR2_X2 U192 ( .A(\eq_169_2/B[4] ), .B(\eq_162_2/A[4] ), .Z(n175) );
  XNOR2_X2 U193 ( .A(\eq_169_2/B[6] ), .B(\eq_162_2/A[6] ), .ZN(n168) );
  XNOR2_X2 U194 ( .A(\eq_169_2/B[7] ), .B(\eq_162_2/A[7] ), .ZN(n167) );
  AND4_X2 U195 ( .A1(n178), .A2(n179), .A3(n180), .A4(n181), .ZN(n155) );
  NOR4_X2 U196 ( .A1(n182), .A2(n183), .A3(n184), .A4(n185), .ZN(n181) );
  XOR2_X2 U197 ( .A(\eq_169_2/B[0] ), .B(\eq_169_2/A[0] ), .Z(n185) );
  XOR2_X2 U198 ( .A(\eq_169_2/B[2] ), .B(\eq_169_2/A[2] ), .Z(n184) );
  XOR2_X2 U199 ( .A(\eq_169_2/B[1] ), .B(\eq_169_2/A[1] ), .Z(n183) );
  NAND3_X2 U200 ( .A1(NewRowY[62]), .A2(NewRowY[61]), .A3(NewRowY[63]), .ZN(
        n182) );
  NOR3_X2 U201 ( .A1(n186), .A2(n187), .A3(n188), .ZN(n180) );
  XOR2_X2 U202 ( .A(\eq_169_2/B[3] ), .B(\eq_169_2/A[3] ), .Z(n188) );
  XOR2_X2 U203 ( .A(\eq_169_2/B[5] ), .B(\eq_169_2/A[5] ), .Z(n187) );
  XOR2_X2 U204 ( .A(\eq_169_2/B[4] ), .B(\eq_169_2/A[4] ), .Z(n186) );
  XNOR2_X2 U205 ( .A(\eq_169_2/B[6] ), .B(\eq_169_2/A[6] ), .ZN(n179) );
  XNOR2_X2 U206 ( .A(\eq_169_2/B[7] ), .B(\eq_169_2/A[7] ), .ZN(n178) );
  NAND4_X2 U207 ( .A1(n189), .A2(n190), .A3(n191), .A4(n192), .ZN(n37) );
  NOR4_X2 U208 ( .A1(n193), .A2(n194), .A3(n195), .A4(n196), .ZN(n192) );
  XOR2_X2 U209 ( .A(\eq_169_2/B[0] ), .B(\eq_147_2/A[0] ), .Z(n196) );
  XOR2_X2 U210 ( .A(\eq_169_2/B[2] ), .B(\eq_147_2/A[2] ), .Z(n195) );
  XOR2_X2 U211 ( .A(\eq_169_2/B[1] ), .B(\eq_147_2/A[1] ), .Z(n194) );
  NAND3_X2 U212 ( .A1(NewRowY[254]), .A2(NewRowY[253]), .A3(NewRowY[255]), 
        .ZN(n193) );
  NOR3_X2 U213 ( .A1(n197), .A2(n198), .A3(n199), .ZN(n191) );
  XOR2_X2 U214 ( .A(\eq_169_2/B[3] ), .B(\eq_147_2/A[3] ), .Z(n199) );
  XOR2_X2 U215 ( .A(\eq_169_2/B[5] ), .B(\eq_147_2/A[5] ), .Z(n198) );
  XOR2_X2 U216 ( .A(\eq_169_2/B[4] ), .B(\eq_147_2/A[4] ), .Z(n197) );
  XNOR2_X2 U217 ( .A(\eq_169_2/B[6] ), .B(\eq_147_2/A[6] ), .ZN(n190) );
  XNOR2_X2 U218 ( .A(\eq_169_2/B[7] ), .B(\eq_147_2/A[7] ), .ZN(n189) );
  NAND2_X2 U220 ( .A1(PosDX[0]), .A2(n900), .ZN(n201) );
  NAND2_X2 U223 ( .A1(PosDX[1]), .A2(n900), .ZN(n206) );
  OAI22_X2 U236 ( .A1(n902), .A2(n901), .B1(n220), .B2(n1), .ZN(n418) );
  NAND2_X2 U237 ( .A1(n221), .A2(n222), .ZN(n419) );
  NAND2_X2 U240 ( .A1(n225), .A2(n226), .ZN(n420) );
  NAND2_X2 U243 ( .A1(n227), .A2(n228), .ZN(n421) );
  NAND2_X2 U246 ( .A1(n229), .A2(n230), .ZN(n422) );
  NAND2_X2 U249 ( .A1(n231), .A2(n232), .ZN(n423) );
  NAND2_X2 U252 ( .A1(n233), .A2(n234), .ZN(n424) );
  NAND2_X2 U255 ( .A1(n235), .A2(n236), .ZN(n425) );
  NAND2_X2 U258 ( .A1(n237), .A2(n238), .ZN(n426) );
  NAND2_X2 U261 ( .A1(n239), .A2(n240), .ZN(n427) );
  NAND2_X2 U264 ( .A1(n241), .A2(n242), .ZN(n428) );
  NAND2_X2 U267 ( .A1(n243), .A2(n244), .ZN(n429) );
  NAND2_X2 U270 ( .A1(n245), .A2(n246), .ZN(n430) );
  NAND2_X2 U273 ( .A1(n247), .A2(n248), .ZN(n431) );
  NAND2_X2 U276 ( .A1(n249), .A2(n250), .ZN(n432) );
  NAND2_X2 U279 ( .A1(n251), .A2(n252), .ZN(n433) );
  NAND2_X2 U282 ( .A1(n253), .A2(n254), .ZN(n434) );
  NAND2_X2 U285 ( .A1(n255), .A2(n256), .ZN(n435) );
  NAND2_X2 U288 ( .A1(n257), .A2(n258), .ZN(n436) );
  NAND2_X2 U291 ( .A1(n259), .A2(n260), .ZN(n437) );
  NAND2_X2 U294 ( .A1(n261), .A2(n262), .ZN(n438) );
  NAND2_X2 U297 ( .A1(n263), .A2(n264), .ZN(n439) );
  NAND2_X2 U300 ( .A1(n265), .A2(n266), .ZN(n440) );
  NAND2_X2 U303 ( .A1(n267), .A2(n268), .ZN(n441) );
  NAND2_X2 U306 ( .A1(n269), .A2(n270), .ZN(n442) );
  NAND2_X2 U309 ( .A1(n271), .A2(n272), .ZN(n443) );
  NAND2_X2 U312 ( .A1(n273), .A2(n274), .ZN(n444) );
  NAND2_X2 U315 ( .A1(n275), .A2(n276), .ZN(n445) );
  NAND2_X2 U318 ( .A1(n277), .A2(n278), .ZN(n446) );
  NAND2_X2 U321 ( .A1(n279), .A2(n280), .ZN(n447) );
  NAND2_X2 U324 ( .A1(n281), .A2(n282), .ZN(n448) );
  NAND2_X2 U327 ( .A1(n283), .A2(n284), .ZN(n449) );
  NAND2_X2 U330 ( .A1(n285), .A2(n286), .ZN(n450) );
  NAND2_X2 U333 ( .A1(n287), .A2(n288), .ZN(n451) );
  NAND2_X2 U336 ( .A1(n289), .A2(n290), .ZN(n452) );
  NAND2_X2 U339 ( .A1(n291), .A2(n292), .ZN(n453) );
  NAND2_X2 U342 ( .A1(n293), .A2(n294), .ZN(n454) );
  NAND2_X2 U345 ( .A1(n295), .A2(n296), .ZN(n455) );
  NAND2_X2 U348 ( .A1(n297), .A2(n298), .ZN(n456) );
  NAND2_X2 U351 ( .A1(n299), .A2(n300), .ZN(n457) );
  NAND2_X2 U354 ( .A1(n301), .A2(n302), .ZN(n458) );
  NAND2_X2 U357 ( .A1(n303), .A2(n304), .ZN(n459) );
  NAND2_X2 U360 ( .A1(n305), .A2(n306), .ZN(n460) );
  NAND2_X2 U363 ( .A1(n307), .A2(n308), .ZN(n461) );
  NAND2_X2 U366 ( .A1(n309), .A2(n310), .ZN(n462) );
  NAND2_X2 U369 ( .A1(n311), .A2(n312), .ZN(n463) );
  NAND2_X2 U372 ( .A1(n313), .A2(n314), .ZN(n464) );
  NAND2_X2 U375 ( .A1(n315), .A2(n316), .ZN(n465) );
  NAND2_X2 U378 ( .A1(n317), .A2(n318), .ZN(n466) );
  NOR2_X2 U380 ( .A1(n202), .A2(n205), .ZN(n224) );
  NAND2_X2 U384 ( .A1(n219), .A2(n154), .ZN(n220) );
  NOR2_X2 U385 ( .A1(EnableChange), .A2(reset), .ZN(n154) );
  NOR3_X2 U386 ( .A1(n320), .A2(n904), .A3(n205), .ZN(n219) );
  NAND2_X2 U387 ( .A1(n319), .A2(n203), .ZN(n205) );
  NAND4_X2 U388 ( .A1(n321), .A2(n322), .A3(n323), .A4(n324), .ZN(n319) );
  NOR4_X2 U389 ( .A1(n325), .A2(n326), .A3(n327), .A4(n328), .ZN(n324) );
  XOR2_X2 U390 ( .A(\eq_63_2/B[0] ), .B(\eq_49_2/A[0] ), .Z(n328) );
  XOR2_X2 U391 ( .A(\eq_63_2/B[2] ), .B(\eq_49_2/A[2] ), .Z(n327) );
  XOR2_X2 U392 ( .A(\eq_63_2/B[1] ), .B(\eq_49_2/A[1] ), .Z(n326) );
  NAND3_X2 U393 ( .A1(NewRowX[190]), .A2(NewRowX[189]), .A3(NewRowX[191]), 
        .ZN(n325) );
  NOR3_X2 U394 ( .A1(n329), .A2(n330), .A3(n331), .ZN(n323) );
  XOR2_X2 U395 ( .A(\eq_63_2/B[3] ), .B(\eq_49_2/A[3] ), .Z(n331) );
  XOR2_X2 U396 ( .A(\eq_63_2/B[5] ), .B(\eq_49_2/A[5] ), .Z(n330) );
  XOR2_X2 U397 ( .A(\eq_63_2/B[4] ), .B(\eq_49_2/A[4] ), .Z(n329) );
  XNOR2_X2 U398 ( .A(\eq_63_2/B[6] ), .B(\eq_49_2/A[6] ), .ZN(n322) );
  XNOR2_X2 U399 ( .A(\eq_63_2/B[7] ), .B(\eq_49_2/A[7] ), .ZN(n321) );
  NAND4_X2 U400 ( .A1(n332), .A2(n333), .A3(n334), .A4(n335), .ZN(n202) );
  NOR4_X2 U401 ( .A1(n336), .A2(n337), .A3(n338), .A4(n339), .ZN(n335) );
  XOR2_X2 U402 ( .A(\eq_63_2/B[0] ), .B(\eq_56_2/A[0] ), .Z(n339) );
  XOR2_X2 U403 ( .A(\eq_63_2/B[2] ), .B(\eq_56_2/A[2] ), .Z(n338) );
  XOR2_X2 U404 ( .A(\eq_63_2/B[1] ), .B(\eq_56_2/A[1] ), .Z(n337) );
  NAND3_X2 U405 ( .A1(NewRowX[126]), .A2(NewRowX[125]), .A3(NewRowX[127]), 
        .ZN(n336) );
  NOR3_X2 U406 ( .A1(n340), .A2(n341), .A3(n342), .ZN(n334) );
  XOR2_X2 U407 ( .A(\eq_63_2/B[3] ), .B(\eq_56_2/A[3] ), .Z(n342) );
  XOR2_X2 U408 ( .A(\eq_63_2/B[5] ), .B(\eq_56_2/A[5] ), .Z(n341) );
  XOR2_X2 U409 ( .A(\eq_63_2/B[4] ), .B(\eq_56_2/A[4] ), .Z(n340) );
  XNOR2_X2 U410 ( .A(\eq_63_2/B[6] ), .B(\eq_56_2/A[6] ), .ZN(n333) );
  XNOR2_X2 U411 ( .A(\eq_63_2/B[7] ), .B(\eq_56_2/A[7] ), .ZN(n332) );
  AND4_X2 U412 ( .A1(n343), .A2(n344), .A3(n345), .A4(n346), .ZN(n320) );
  NOR4_X2 U413 ( .A1(n347), .A2(n348), .A3(n349), .A4(n350), .ZN(n346) );
  XOR2_X2 U414 ( .A(\eq_63_2/B[0] ), .B(\eq_63_2/A[0] ), .Z(n350) );
  XOR2_X2 U415 ( .A(\eq_63_2/B[2] ), .B(\eq_63_2/A[2] ), .Z(n349) );
  XOR2_X2 U416 ( .A(\eq_63_2/B[1] ), .B(\eq_63_2/A[1] ), .Z(n348) );
  NAND3_X2 U417 ( .A1(NewRowX[62]), .A2(NewRowX[61]), .A3(NewRowX[63]), .ZN(
        n347) );
  NOR3_X2 U418 ( .A1(n351), .A2(n352), .A3(n353), .ZN(n345) );
  XOR2_X2 U419 ( .A(\eq_63_2/B[3] ), .B(\eq_63_2/A[3] ), .Z(n353) );
  XOR2_X2 U420 ( .A(\eq_63_2/B[5] ), .B(\eq_63_2/A[5] ), .Z(n352) );
  XOR2_X2 U421 ( .A(\eq_63_2/B[4] ), .B(\eq_63_2/A[4] ), .Z(n351) );
  XNOR2_X2 U422 ( .A(\eq_63_2/B[6] ), .B(\eq_63_2/A[6] ), .ZN(n344) );
  XNOR2_X2 U423 ( .A(\eq_63_2/B[7] ), .B(\eq_63_2/A[7] ), .ZN(n343) );
  NAND4_X2 U424 ( .A1(n354), .A2(n355), .A3(n356), .A4(n357), .ZN(n203) );
  NOR4_X2 U425 ( .A1(n358), .A2(n359), .A3(n360), .A4(n361), .ZN(n357) );
  XOR2_X2 U426 ( .A(\eq_63_2/B[0] ), .B(\eq_41_2/A[0] ), .Z(n361) );
  XOR2_X2 U427 ( .A(\eq_63_2/B[2] ), .B(\eq_41_2/A[2] ), .Z(n360) );
  XOR2_X2 U428 ( .A(\eq_63_2/B[1] ), .B(\eq_41_2/A[1] ), .Z(n359) );
  NAND3_X2 U429 ( .A1(NewRowX[254]), .A2(NewRowX[253]), .A3(NewRowX[255]), 
        .ZN(n358) );
  NOR3_X2 U430 ( .A1(n362), .A2(n363), .A3(n364), .ZN(n356) );
  XOR2_X2 U431 ( .A(\eq_63_2/B[3] ), .B(\eq_41_2/A[3] ), .Z(n364) );
  XOR2_X2 U432 ( .A(\eq_63_2/B[5] ), .B(\eq_41_2/A[5] ), .Z(n363) );
  XOR2_X2 U433 ( .A(\eq_63_2/B[4] ), .B(\eq_41_2/A[4] ), .Z(n362) );
  XNOR2_X2 U434 ( .A(\eq_63_2/B[6] ), .B(\eq_41_2/A[6] ), .ZN(n355) );
  XNOR2_X2 U435 ( .A(\eq_63_2/B[7] ), .B(\eq_41_2/A[7] ), .ZN(n354) );
  DFF_X2 DiagonalDoneY_reg ( .D(n367), .CK(clock), .Q(DiagonalDoneY), .QN(n13)
         );
  DFF_X2 DiagonalDoneX_reg ( .D(n418), .CK(clock), .Q(DiagonalDoneX), .QN(n1)
         );
  NOR3_X4 U3 ( .A1(n903), .A2(n906), .A3(n39), .ZN(n867) );
  NOR2_X4 U5 ( .A1(n319), .A2(n872), .ZN(n868) );
  NOR2_X4 U6 ( .A1(n153), .A2(n905), .ZN(n869) );
  NOR2_X4 U8 ( .A1(n36), .A2(n39), .ZN(n870) );
  OR3_X4 U9 ( .A1(n902), .A2(n904), .A3(n205), .ZN(n871) );
  INV_X4 U10 ( .A(n871), .ZN(n876) );
  INV_X4 U11 ( .A(n871), .ZN(n875) );
  INV_X4 U12 ( .A(n874), .ZN(n873) );
  INV_X4 U13 ( .A(n203), .ZN(n872) );
  INV_X4 U14 ( .A(n42), .ZN(n899) );
  INV_X4 U15 ( .A(n208), .ZN(n900) );
  INV_X4 U16 ( .A(n224), .ZN(n874) );
  NOR2_X2 U17 ( .A1(n901), .A2(n53), .ZN(n42) );
  NOR2_X2 U18 ( .A1(n901), .A2(n219), .ZN(n208) );
  AOI22_X2 U19 ( .A1(\U3/U10/DATA1_0 ), .A2(n872), .B1(DiagonalX[0]), .B2(n902), .ZN(n221) );
  AOI222_X1 U22 ( .A1(\U3/U10/DATA2_0 ), .A2(n868), .B1(\U3/U10/DATA4_0 ), 
        .B2(n876), .C1(\U3/U10/DATA3_0 ), .C2(n873), .ZN(n222) );
  AOI22_X2 U23 ( .A1(\U3/U10/DATA1_1 ), .A2(n872), .B1(DiagonalX[1]), .B2(n902), .ZN(n225) );
  AOI222_X1 U25 ( .A1(\U3/U10/DATA2_1 ), .A2(n868), .B1(\U3/U10/DATA4_1 ), 
        .B2(n876), .C1(\U3/U10/DATA3_1 ), .C2(n873), .ZN(n226) );
  AOI22_X2 U26 ( .A1(\U3/U10/DATA1_2 ), .A2(n872), .B1(DiagonalX[2]), .B2(n902), .ZN(n227) );
  AOI222_X1 U28 ( .A1(\U3/U10/DATA2_2 ), .A2(n868), .B1(\U3/U10/DATA4_2 ), 
        .B2(n876), .C1(\U3/U10/DATA3_2 ), .C2(n873), .ZN(n228) );
  AOI22_X2 U29 ( .A1(\U3/U10/DATA1_3 ), .A2(n872), .B1(DiagonalX[3]), .B2(n902), .ZN(n229) );
  AOI222_X1 U31 ( .A1(\U3/U10/DATA2_3 ), .A2(n868), .B1(\U3/U10/DATA4_3 ), 
        .B2(n876), .C1(\U3/U10/DATA3_3 ), .C2(n873), .ZN(n230) );
  AOI22_X2 U32 ( .A1(\U3/U10/DATA1_4 ), .A2(n872), .B1(DiagonalX[4]), .B2(n902), .ZN(n231) );
  AOI222_X1 U34 ( .A1(\U3/U10/DATA2_4 ), .A2(n868), .B1(\U3/U10/DATA4_4 ), 
        .B2(n876), .C1(\U3/U10/DATA3_4 ), .C2(n873), .ZN(n232) );
  AOI22_X2 U35 ( .A1(\U3/U10/DATA1_5 ), .A2(n872), .B1(DiagonalX[5]), .B2(n902), .ZN(n233) );
  AOI222_X1 U37 ( .A1(\U3/U10/DATA2_5 ), .A2(n868), .B1(\U3/U10/DATA4_5 ), 
        .B2(n876), .C1(\U3/U10/DATA3_5 ), .C2(n873), .ZN(n234) );
  AOI22_X2 U38 ( .A1(\U3/U10/DATA1_6 ), .A2(n872), .B1(DiagonalX[6]), .B2(n902), .ZN(n235) );
  AOI222_X1 U40 ( .A1(\U3/U10/DATA2_6 ), .A2(n868), .B1(\U3/U10/DATA4_6 ), 
        .B2(n876), .C1(\U3/U10/DATA3_6 ), .C2(n873), .ZN(n236) );
  AOI22_X2 U41 ( .A1(\U3/U10/DATA1_7 ), .A2(n872), .B1(DiagonalX[7]), .B2(n902), .ZN(n237) );
  AOI222_X1 U43 ( .A1(\U3/U10/DATA2_7 ), .A2(n868), .B1(\U3/U10/DATA4_7 ), 
        .B2(n876), .C1(\U3/U10/DATA3_7 ), .C2(n873), .ZN(n238) );
  AOI22_X2 U44 ( .A1(\U3/U10/DATA1_8 ), .A2(n872), .B1(DiagonalX[8]), .B2(n902), .ZN(n239) );
  AOI222_X1 U46 ( .A1(\U3/U10/DATA2_8 ), .A2(n868), .B1(\U3/U10/DATA4_8 ), 
        .B2(n876), .C1(\U3/U10/DATA3_8 ), .C2(n873), .ZN(n240) );
  AOI22_X2 U47 ( .A1(\U3/U10/DATA1_9 ), .A2(n872), .B1(DiagonalX[9]), .B2(n902), .ZN(n241) );
  AOI222_X1 U49 ( .A1(\U3/U10/DATA2_9 ), .A2(n868), .B1(\U3/U10/DATA4_9 ), 
        .B2(n876), .C1(\U3/U10/DATA3_9 ), .C2(n873), .ZN(n242) );
  AOI22_X2 U50 ( .A1(\U3/U10/DATA1_10 ), .A2(n872), .B1(DiagonalX[10]), .B2(
        n902), .ZN(n243) );
  AOI222_X1 U52 ( .A1(\U3/U10/DATA2_10 ), .A2(n868), .B1(\U3/U10/DATA4_10 ), 
        .B2(n876), .C1(\U3/U10/DATA3_10 ), .C2(n873), .ZN(n244) );
  AOI22_X2 U53 ( .A1(\U3/U10/DATA1_11 ), .A2(n872), .B1(DiagonalX[11]), .B2(
        n902), .ZN(n245) );
  AOI222_X1 U55 ( .A1(\U3/U10/DATA2_11 ), .A2(n868), .B1(\U3/U10/DATA4_11 ), 
        .B2(n876), .C1(\U3/U10/DATA3_11 ), .C2(n873), .ZN(n246) );
  AOI22_X2 U56 ( .A1(\U3/U10/DATA1_12 ), .A2(n872), .B1(DiagonalX[12]), .B2(
        n902), .ZN(n247) );
  AOI222_X1 U58 ( .A1(\U3/U10/DATA2_12 ), .A2(n868), .B1(\U3/U10/DATA4_12 ), 
        .B2(n875), .C1(\U3/U10/DATA3_12 ), .C2(n224), .ZN(n248) );
  AOI22_X2 U59 ( .A1(\U3/U10/DATA1_13 ), .A2(n872), .B1(DiagonalX[13]), .B2(
        n902), .ZN(n249) );
  AOI222_X1 U61 ( .A1(\U3/U10/DATA2_13 ), .A2(n868), .B1(\U3/U10/DATA4_13 ), 
        .B2(n875), .C1(\U3/U10/DATA3_13 ), .C2(n224), .ZN(n250) );
  AOI22_X2 U62 ( .A1(\U3/U10/DATA1_14 ), .A2(n872), .B1(DiagonalX[14]), .B2(
        n902), .ZN(n251) );
  AOI222_X1 U64 ( .A1(\U3/U10/DATA2_14 ), .A2(n868), .B1(\U3/U10/DATA4_14 ), 
        .B2(n875), .C1(\U3/U10/DATA3_14 ), .C2(n224), .ZN(n252) );
  AOI22_X2 U65 ( .A1(\U3/U10/DATA1_15 ), .A2(n872), .B1(DiagonalX[15]), .B2(
        n902), .ZN(n253) );
  AOI222_X1 U67 ( .A1(\U3/U10/DATA2_15 ), .A2(n868), .B1(\U3/U10/DATA4_15 ), 
        .B2(n875), .C1(\U3/U10/DATA3_15 ), .C2(n224), .ZN(n254) );
  AOI22_X2 U68 ( .A1(\U3/U10/DATA1_16 ), .A2(n872), .B1(DiagonalX[16]), .B2(
        n902), .ZN(n255) );
  AOI222_X1 U70 ( .A1(\U3/U10/DATA2_16 ), .A2(n868), .B1(\U3/U10/DATA4_16 ), 
        .B2(n875), .C1(\U3/U10/DATA3_16 ), .C2(n224), .ZN(n256) );
  AOI22_X2 U71 ( .A1(\U3/U10/DATA1_17 ), .A2(n872), .B1(DiagonalX[17]), .B2(
        n902), .ZN(n257) );
  AOI222_X1 U73 ( .A1(\U3/U10/DATA2_17 ), .A2(n868), .B1(\U3/U10/DATA4_17 ), 
        .B2(n875), .C1(\U3/U10/DATA3_17 ), .C2(n224), .ZN(n258) );
  AOI22_X2 U74 ( .A1(\U3/U10/DATA1_18 ), .A2(n872), .B1(DiagonalX[18]), .B2(
        n902), .ZN(n259) );
  AOI222_X1 U76 ( .A1(\U3/U10/DATA2_18 ), .A2(n868), .B1(\U3/U10/DATA4_18 ), 
        .B2(n875), .C1(\U3/U10/DATA3_18 ), .C2(n224), .ZN(n260) );
  AOI22_X2 U77 ( .A1(\U3/U10/DATA1_19 ), .A2(n872), .B1(DiagonalX[19]), .B2(
        n902), .ZN(n261) );
  AOI222_X1 U79 ( .A1(\U3/U10/DATA2_19 ), .A2(n868), .B1(\U3/U10/DATA4_19 ), 
        .B2(n875), .C1(\U3/U10/DATA3_19 ), .C2(n224), .ZN(n262) );
  AOI22_X2 U80 ( .A1(\U3/U10/DATA1_20 ), .A2(n872), .B1(DiagonalX[20]), .B2(
        n902), .ZN(n263) );
  AOI222_X1 U82 ( .A1(\U3/U10/DATA2_20 ), .A2(n868), .B1(\U3/U10/DATA4_20 ), 
        .B2(n875), .C1(\U3/U10/DATA3_20 ), .C2(n224), .ZN(n264) );
  AOI22_X2 U83 ( .A1(\U3/U10/DATA1_21 ), .A2(n872), .B1(DiagonalX[21]), .B2(
        n902), .ZN(n265) );
  AOI222_X1 U85 ( .A1(\U3/U10/DATA2_21 ), .A2(n868), .B1(\U3/U10/DATA4_21 ), 
        .B2(n875), .C1(\U3/U10/DATA3_21 ), .C2(n224), .ZN(n266) );
  AOI22_X2 U86 ( .A1(\U3/U10/DATA1_22 ), .A2(n872), .B1(DiagonalX[22]), .B2(
        n902), .ZN(n267) );
  AOI222_X1 U88 ( .A1(\U3/U10/DATA2_22 ), .A2(n868), .B1(\U3/U10/DATA4_22 ), 
        .B2(n875), .C1(\U3/U10/DATA3_22 ), .C2(n224), .ZN(n268) );
  AOI22_X2 U89 ( .A1(\U3/U10/DATA1_23 ), .A2(n872), .B1(DiagonalX[23]), .B2(
        n902), .ZN(n269) );
  AOI222_X1 U91 ( .A1(\U3/U10/DATA2_23 ), .A2(n868), .B1(\U3/U10/DATA4_23 ), 
        .B2(n875), .C1(\U3/U10/DATA3_23 ), .C2(n224), .ZN(n270) );
  AOI22_X2 U92 ( .A1(\U3/U10/DATA1_24 ), .A2(n872), .B1(DiagonalX[24]), .B2(
        n902), .ZN(n271) );
  AOI222_X1 U94 ( .A1(\U3/U10/DATA2_24 ), .A2(n868), .B1(\U3/U10/DATA4_24 ), 
        .B2(n876), .C1(\U3/U10/DATA3_24 ), .C2(n873), .ZN(n272) );
  AOI22_X2 U95 ( .A1(\U3/U10/DATA1_25 ), .A2(n872), .B1(DiagonalX[25]), .B2(
        n902), .ZN(n273) );
  AOI222_X1 U97 ( .A1(\U3/U10/DATA2_25 ), .A2(n868), .B1(\U3/U10/DATA4_25 ), 
        .B2(n875), .C1(\U3/U10/DATA3_25 ), .C2(n873), .ZN(n274) );
  AOI22_X2 U98 ( .A1(\U3/U10/DATA1_26 ), .A2(n872), .B1(DiagonalX[26]), .B2(
        n902), .ZN(n275) );
  AOI222_X1 U100 ( .A1(\U3/U10/DATA2_26 ), .A2(n868), .B1(\U3/U10/DATA4_26 ), 
        .B2(n876), .C1(\U3/U10/DATA3_26 ), .C2(n873), .ZN(n276) );
  AOI22_X2 U101 ( .A1(\U3/U10/DATA1_27 ), .A2(n872), .B1(DiagonalX[27]), .B2(
        n902), .ZN(n277) );
  AOI222_X1 U103 ( .A1(\U3/U10/DATA2_27 ), .A2(n868), .B1(\U3/U10/DATA4_27 ), 
        .B2(n875), .C1(\U3/U10/DATA3_27 ), .C2(n224), .ZN(n278) );
  AOI22_X2 U104 ( .A1(\U3/U10/DATA1_28 ), .A2(n872), .B1(DiagonalX[28]), .B2(
        n902), .ZN(n279) );
  AOI222_X1 U106 ( .A1(\U3/U10/DATA2_28 ), .A2(n868), .B1(\U3/U10/DATA4_28 ), 
        .B2(n876), .C1(\U3/U10/DATA3_28 ), .C2(n224), .ZN(n280) );
  AOI22_X2 U107 ( .A1(\U3/U10/DATA1_29 ), .A2(n872), .B1(DiagonalX[29]), .B2(
        n902), .ZN(n281) );
  AOI222_X1 U109 ( .A1(\U3/U10/DATA2_29 ), .A2(n868), .B1(\U3/U10/DATA4_29 ), 
        .B2(n875), .C1(\U3/U10/DATA3_29 ), .C2(n224), .ZN(n282) );
  AOI22_X2 U110 ( .A1(\U3/U10/DATA1_30 ), .A2(n872), .B1(DiagonalX[30]), .B2(
        n902), .ZN(n283) );
  AOI222_X1 U112 ( .A1(\U3/U10/DATA2_30 ), .A2(n868), .B1(\U3/U10/DATA4_30 ), 
        .B2(n876), .C1(\U3/U10/DATA3_30 ), .C2(n224), .ZN(n284) );
  AOI22_X2 U113 ( .A1(\U3/U10/DATA1_31 ), .A2(n872), .B1(DiagonalX[31]), .B2(
        n902), .ZN(n285) );
  AOI222_X1 U115 ( .A1(\U3/U10/DATA2_31 ), .A2(n868), .B1(\U3/U10/DATA4_31 ), 
        .B2(n875), .C1(\U3/U10/DATA3_31 ), .C2(n224), .ZN(n286) );
  AOI22_X2 U116 ( .A1(\U3/U10/DATA1_32 ), .A2(n872), .B1(DiagonalX[32]), .B2(
        n902), .ZN(n287) );
  AOI222_X1 U118 ( .A1(\U3/U10/DATA2_32 ), .A2(n868), .B1(\U3/U10/DATA4_32 ), 
        .B2(n876), .C1(\U3/U10/DATA3_32 ), .C2(n224), .ZN(n288) );
  AOI22_X2 U119 ( .A1(\U3/U10/DATA1_33 ), .A2(n872), .B1(DiagonalX[33]), .B2(
        n902), .ZN(n289) );
  AOI222_X1 U121 ( .A1(\U3/U10/DATA2_33 ), .A2(n868), .B1(\U3/U10/DATA4_33 ), 
        .B2(n875), .C1(\U3/U10/DATA3_33 ), .C2(n224), .ZN(n290) );
  AOI22_X2 U122 ( .A1(\U3/U10/DATA1_34 ), .A2(n872), .B1(DiagonalX[34]), .B2(
        n902), .ZN(n291) );
  AOI222_X1 U124 ( .A1(\U3/U10/DATA2_34 ), .A2(n868), .B1(\U3/U10/DATA4_34 ), 
        .B2(n876), .C1(\U3/U10/DATA3_34 ), .C2(n224), .ZN(n292) );
  AOI22_X2 U125 ( .A1(\U3/U10/DATA1_35 ), .A2(n872), .B1(DiagonalX[35]), .B2(
        n902), .ZN(n293) );
  AOI222_X1 U127 ( .A1(\U3/U10/DATA2_35 ), .A2(n868), .B1(\U3/U10/DATA4_35 ), 
        .B2(n875), .C1(\U3/U10/DATA3_35 ), .C2(n224), .ZN(n294) );
  AOI22_X2 U128 ( .A1(\U3/U10/DATA1_36 ), .A2(n872), .B1(DiagonalX[36]), .B2(
        n902), .ZN(n295) );
  AOI222_X1 U130 ( .A1(\U3/U10/DATA2_36 ), .A2(n868), .B1(\U3/U10/DATA4_36 ), 
        .B2(n876), .C1(\U3/U10/DATA3_36 ), .C2(n873), .ZN(n296) );
  AOI22_X2 U131 ( .A1(\U3/U10/DATA1_37 ), .A2(n872), .B1(DiagonalX[37]), .B2(
        n902), .ZN(n297) );
  AOI222_X1 U133 ( .A1(\U3/U10/DATA2_37 ), .A2(n868), .B1(\U3/U10/DATA4_37 ), 
        .B2(n876), .C1(\U3/U10/DATA3_37 ), .C2(n224), .ZN(n298) );
  AOI22_X2 U134 ( .A1(\U3/U10/DATA1_38 ), .A2(n872), .B1(DiagonalX[38]), .B2(
        n902), .ZN(n299) );
  AOI222_X1 U136 ( .A1(\U3/U10/DATA2_38 ), .A2(n868), .B1(\U3/U10/DATA4_38 ), 
        .B2(n875), .C1(\U3/U10/DATA3_38 ), .C2(n873), .ZN(n300) );
  AOI22_X2 U137 ( .A1(\U3/U10/DATA1_39 ), .A2(n872), .B1(DiagonalX[39]), .B2(
        n902), .ZN(n301) );
  AOI222_X1 U139 ( .A1(\U3/U10/DATA2_39 ), .A2(n868), .B1(\U3/U10/DATA4_39 ), 
        .B2(n875), .C1(\U3/U10/DATA3_39 ), .C2(n224), .ZN(n302) );
  AOI22_X2 U140 ( .A1(\U3/U10/DATA1_40 ), .A2(n872), .B1(DiagonalX[40]), .B2(
        n902), .ZN(n303) );
  AOI222_X1 U142 ( .A1(\U3/U10/DATA2_40 ), .A2(n868), .B1(\U3/U10/DATA4_40 ), 
        .B2(n876), .C1(\U3/U10/DATA3_40 ), .C2(n224), .ZN(n304) );
  AOI22_X2 U143 ( .A1(\U3/U10/DATA1_41 ), .A2(n872), .B1(DiagonalX[41]), .B2(
        n902), .ZN(n305) );
  AOI222_X1 U145 ( .A1(\U3/U10/DATA2_41 ), .A2(n868), .B1(\U3/U10/DATA4_41 ), 
        .B2(n875), .C1(\U3/U10/DATA3_41 ), .C2(n224), .ZN(n306) );
  AOI22_X2 U146 ( .A1(\U3/U10/DATA1_42 ), .A2(n872), .B1(DiagonalX[42]), .B2(
        n902), .ZN(n307) );
  AOI222_X1 U148 ( .A1(\U3/U10/DATA2_42 ), .A2(n868), .B1(\U3/U10/DATA4_42 ), 
        .B2(n876), .C1(\U3/U10/DATA3_42 ), .C2(n224), .ZN(n308) );
  AOI22_X2 U149 ( .A1(\U3/U10/DATA1_43 ), .A2(n872), .B1(DiagonalX[43]), .B2(
        n902), .ZN(n309) );
  AOI222_X1 U151 ( .A1(\U3/U10/DATA2_43 ), .A2(n868), .B1(\U3/U10/DATA4_43 ), 
        .B2(n876), .C1(\U3/U10/DATA3_43 ), .C2(n224), .ZN(n310) );
  AOI22_X2 U152 ( .A1(\U3/U10/DATA1_44 ), .A2(n872), .B1(DiagonalX[44]), .B2(
        n902), .ZN(n311) );
  AOI222_X1 U154 ( .A1(\U3/U10/DATA2_44 ), .A2(n868), .B1(\U3/U10/DATA4_44 ), 
        .B2(n875), .C1(\U3/U10/DATA3_44 ), .C2(n224), .ZN(n312) );
  AOI22_X2 U155 ( .A1(\U3/U10/DATA1_45 ), .A2(n872), .B1(DiagonalX[45]), .B2(
        n902), .ZN(n313) );
  AOI222_X1 U157 ( .A1(\U3/U10/DATA2_45 ), .A2(n868), .B1(\U3/U10/DATA4_45 ), 
        .B2(n875), .C1(\U3/U10/DATA3_45 ), .C2(n224), .ZN(n314) );
  AOI22_X2 U158 ( .A1(\U3/U10/DATA1_46 ), .A2(n872), .B1(DiagonalX[46]), .B2(
        n902), .ZN(n315) );
  AOI222_X1 U160 ( .A1(\U3/U10/DATA2_46 ), .A2(n868), .B1(\U3/U10/DATA4_46 ), 
        .B2(n876), .C1(\U3/U10/DATA3_46 ), .C2(n224), .ZN(n316) );
  AOI22_X2 U161 ( .A1(\U3/U10/DATA1_47 ), .A2(n872), .B1(DiagonalX[47]), .B2(
        n902), .ZN(n317) );
  AOI222_X1 U163 ( .A1(\U3/U10/DATA2_47 ), .A2(n868), .B1(\U3/U10/DATA4_47 ), 
        .B2(n875), .C1(\U3/U10/DATA3_47 ), .C2(n224), .ZN(n318) );
  AOI22_X2 U164 ( .A1(PosDY[2]), .A2(n899), .B1(Row_noY[0]), .B2(n42), .ZN(n41) );
  AOI22_X2 U165 ( .A1(PosDY[3]), .A2(n899), .B1(Row_noY[1]), .B2(n42), .ZN(n43) );
  AOI22_X2 U166 ( .A1(PosDY[4]), .A2(n899), .B1(Row_noY[2]), .B2(n42), .ZN(n44) );
  AOI22_X2 U167 ( .A1(PosDY[5]), .A2(n899), .B1(Row_noY[3]), .B2(n42), .ZN(n45) );
  AOI22_X2 U219 ( .A1(PosDY[6]), .A2(n899), .B1(Row_noY[4]), .B2(n42), .ZN(n46) );
  AOI22_X2 U221 ( .A1(PosDY[7]), .A2(n899), .B1(Row_noY[5]), .B2(n42), .ZN(n47) );
  AOI22_X2 U222 ( .A1(PosDY[8]), .A2(n899), .B1(Row_noY[6]), .B2(n42), .ZN(n48) );
  AOI22_X2 U224 ( .A1(PosDY[9]), .A2(n899), .B1(Row_noY[7]), .B2(n42), .ZN(n49) );
  AOI22_X2 U225 ( .A1(PosDY[10]), .A2(n899), .B1(Row_noY[8]), .B2(n42), .ZN(
        n50) );
  AOI22_X2 U226 ( .A1(PosDY[11]), .A2(n899), .B1(Row_noY[9]), .B2(n42), .ZN(
        n51) );
  AOI22_X2 U227 ( .A1(PosDY[12]), .A2(n899), .B1(Row_noY[10]), .B2(n42), .ZN(
        n52) );
  OAI21_X2 U228 ( .B1(n200), .B2(n900), .A(n201), .ZN(n416) );
  AOI21_X2 U229 ( .B1(n202), .B2(n203), .A(n868), .ZN(n200) );
  OAI21_X2 U230 ( .B1(n34), .B2(n899), .A(n35), .ZN(n365) );
  AOI21_X2 U231 ( .B1(n36), .B2(n37), .A(n869), .ZN(n34) );
  OAI21_X2 U232 ( .B1(n205), .B2(n900), .A(n206), .ZN(n417) );
  OAI21_X2 U233 ( .B1(n39), .B2(n899), .A(n40), .ZN(n366) );
  AOI22_X2 U234 ( .A1(\U3/U12/DATA1_0 ), .A2(n905), .B1(DiagonalY[0]), .B2(
        n903), .ZN(n55) );
  AOI222_X1 U235 ( .A1(\U3/U12/DATA2_0 ), .A2(n869), .B1(\U3/U12/DATA4_0 ), 
        .B2(n867), .C1(\U3/U12/DATA3_0 ), .C2(n870), .ZN(n56) );
  AOI22_X2 U238 ( .A1(\U3/U12/DATA1_1 ), .A2(n905), .B1(DiagonalY[1]), .B2(
        n903), .ZN(n59) );
  AOI222_X1 U239 ( .A1(\U3/U12/DATA2_1 ), .A2(n869), .B1(\U3/U12/DATA4_1 ), 
        .B2(n867), .C1(\U3/U12/DATA3_1 ), .C2(n870), .ZN(n60) );
  AOI22_X2 U241 ( .A1(\U3/U12/DATA1_2 ), .A2(n905), .B1(DiagonalY[2]), .B2(
        n903), .ZN(n61) );
  AOI222_X1 U242 ( .A1(\U3/U12/DATA2_2 ), .A2(n869), .B1(\U3/U12/DATA4_2 ), 
        .B2(n867), .C1(\U3/U12/DATA3_2 ), .C2(n870), .ZN(n62) );
  AOI22_X2 U244 ( .A1(\U3/U12/DATA1_3 ), .A2(n905), .B1(DiagonalY[3]), .B2(
        n903), .ZN(n63) );
  AOI222_X1 U245 ( .A1(\U3/U12/DATA2_3 ), .A2(n869), .B1(\U3/U12/DATA4_3 ), 
        .B2(n867), .C1(\U3/U12/DATA3_3 ), .C2(n870), .ZN(n64) );
  AOI22_X2 U247 ( .A1(\U3/U12/DATA1_4 ), .A2(n905), .B1(DiagonalY[4]), .B2(
        n903), .ZN(n65) );
  AOI222_X1 U248 ( .A1(\U3/U12/DATA2_4 ), .A2(n869), .B1(\U3/U12/DATA4_4 ), 
        .B2(n867), .C1(\U3/U12/DATA3_4 ), .C2(n870), .ZN(n66) );
  AOI22_X2 U250 ( .A1(\U3/U12/DATA1_5 ), .A2(n905), .B1(DiagonalY[5]), .B2(
        n903), .ZN(n67) );
  AOI222_X1 U251 ( .A1(\U3/U12/DATA2_5 ), .A2(n869), .B1(\U3/U12/DATA4_5 ), 
        .B2(n867), .C1(\U3/U12/DATA3_5 ), .C2(n870), .ZN(n68) );
  AOI22_X2 U253 ( .A1(\U3/U12/DATA1_6 ), .A2(n905), .B1(DiagonalY[6]), .B2(
        n903), .ZN(n69) );
  AOI222_X1 U254 ( .A1(\U3/U12/DATA2_6 ), .A2(n869), .B1(\U3/U12/DATA4_6 ), 
        .B2(n867), .C1(\U3/U12/DATA3_6 ), .C2(n870), .ZN(n70) );
  AOI22_X2 U256 ( .A1(\U3/U12/DATA1_7 ), .A2(n905), .B1(DiagonalY[7]), .B2(
        n903), .ZN(n71) );
  AOI222_X1 U257 ( .A1(\U3/U12/DATA2_7 ), .A2(n869), .B1(\U3/U12/DATA4_7 ), 
        .B2(n867), .C1(\U3/U12/DATA3_7 ), .C2(n870), .ZN(n72) );
  AOI22_X2 U259 ( .A1(\U3/U12/DATA1_8 ), .A2(n905), .B1(DiagonalY[8]), .B2(
        n903), .ZN(n73) );
  AOI222_X1 U260 ( .A1(\U3/U12/DATA2_8 ), .A2(n869), .B1(\U3/U12/DATA4_8 ), 
        .B2(n867), .C1(\U3/U12/DATA3_8 ), .C2(n870), .ZN(n74) );
  AOI22_X2 U262 ( .A1(\U3/U12/DATA1_9 ), .A2(n905), .B1(DiagonalY[9]), .B2(
        n903), .ZN(n75) );
  AOI222_X1 U263 ( .A1(\U3/U12/DATA2_9 ), .A2(n869), .B1(\U3/U12/DATA4_9 ), 
        .B2(n867), .C1(\U3/U12/DATA3_9 ), .C2(n870), .ZN(n76) );
  AOI22_X2 U265 ( .A1(\U3/U12/DATA1_10 ), .A2(n905), .B1(DiagonalY[10]), .B2(
        n903), .ZN(n77) );
  AOI222_X1 U266 ( .A1(\U3/U12/DATA2_10 ), .A2(n869), .B1(\U3/U12/DATA4_10 ), 
        .B2(n867), .C1(\U3/U12/DATA3_10 ), .C2(n870), .ZN(n78) );
  AOI22_X2 U268 ( .A1(\U3/U12/DATA1_11 ), .A2(n905), .B1(DiagonalY[11]), .B2(
        n903), .ZN(n79) );
  AOI222_X1 U269 ( .A1(\U3/U12/DATA2_11 ), .A2(n869), .B1(\U3/U12/DATA4_11 ), 
        .B2(n867), .C1(\U3/U12/DATA3_11 ), .C2(n870), .ZN(n80) );
  AOI22_X2 U271 ( .A1(\U3/U12/DATA1_12 ), .A2(n905), .B1(DiagonalY[12]), .B2(
        n903), .ZN(n81) );
  AOI222_X1 U272 ( .A1(\U3/U12/DATA2_12 ), .A2(n869), .B1(\U3/U12/DATA4_12 ), 
        .B2(n867), .C1(\U3/U12/DATA3_12 ), .C2(n870), .ZN(n82) );
  AOI22_X2 U274 ( .A1(\U3/U12/DATA1_13 ), .A2(n905), .B1(DiagonalY[13]), .B2(
        n903), .ZN(n83) );
  AOI222_X1 U275 ( .A1(\U3/U12/DATA2_13 ), .A2(n869), .B1(\U3/U12/DATA4_13 ), 
        .B2(n867), .C1(\U3/U12/DATA3_13 ), .C2(n870), .ZN(n84) );
  AOI22_X2 U277 ( .A1(\U3/U12/DATA1_14 ), .A2(n905), .B1(DiagonalY[14]), .B2(
        n903), .ZN(n85) );
  AOI222_X1 U278 ( .A1(\U3/U12/DATA2_14 ), .A2(n869), .B1(\U3/U12/DATA4_14 ), 
        .B2(n867), .C1(\U3/U12/DATA3_14 ), .C2(n870), .ZN(n86) );
  AOI22_X2 U280 ( .A1(\U3/U12/DATA1_15 ), .A2(n905), .B1(DiagonalY[15]), .B2(
        n903), .ZN(n87) );
  AOI222_X1 U281 ( .A1(\U3/U12/DATA2_15 ), .A2(n869), .B1(\U3/U12/DATA4_15 ), 
        .B2(n867), .C1(\U3/U12/DATA3_15 ), .C2(n870), .ZN(n88) );
  AOI22_X2 U283 ( .A1(\U3/U12/DATA1_16 ), .A2(n905), .B1(DiagonalY[16]), .B2(
        n903), .ZN(n89) );
  AOI222_X1 U284 ( .A1(\U3/U12/DATA2_16 ), .A2(n869), .B1(\U3/U12/DATA4_16 ), 
        .B2(n867), .C1(\U3/U12/DATA3_16 ), .C2(n870), .ZN(n90) );
  AOI22_X2 U286 ( .A1(\U3/U12/DATA1_17 ), .A2(n905), .B1(DiagonalY[17]), .B2(
        n903), .ZN(n91) );
  AOI222_X1 U287 ( .A1(\U3/U12/DATA2_17 ), .A2(n869), .B1(\U3/U12/DATA4_17 ), 
        .B2(n867), .C1(\U3/U12/DATA3_17 ), .C2(n870), .ZN(n92) );
  AOI22_X2 U289 ( .A1(\U3/U12/DATA1_18 ), .A2(n905), .B1(DiagonalY[18]), .B2(
        n903), .ZN(n93) );
  AOI222_X1 U290 ( .A1(\U3/U12/DATA2_18 ), .A2(n869), .B1(\U3/U12/DATA4_18 ), 
        .B2(n867), .C1(\U3/U12/DATA3_18 ), .C2(n870), .ZN(n94) );
  AOI22_X2 U292 ( .A1(\U3/U12/DATA1_19 ), .A2(n905), .B1(DiagonalY[19]), .B2(
        n903), .ZN(n95) );
  AOI222_X1 U293 ( .A1(\U3/U12/DATA2_19 ), .A2(n869), .B1(\U3/U12/DATA4_19 ), 
        .B2(n867), .C1(\U3/U12/DATA3_19 ), .C2(n870), .ZN(n96) );
  AOI22_X2 U295 ( .A1(\U3/U12/DATA1_20 ), .A2(n905), .B1(DiagonalY[20]), .B2(
        n903), .ZN(n97) );
  AOI222_X1 U296 ( .A1(\U3/U12/DATA2_20 ), .A2(n869), .B1(\U3/U12/DATA4_20 ), 
        .B2(n867), .C1(\U3/U12/DATA3_20 ), .C2(n870), .ZN(n98) );
  AOI22_X2 U298 ( .A1(\U3/U12/DATA1_21 ), .A2(n905), .B1(DiagonalY[21]), .B2(
        n903), .ZN(n99) );
  AOI222_X1 U299 ( .A1(\U3/U12/DATA2_21 ), .A2(n869), .B1(\U3/U12/DATA4_21 ), 
        .B2(n867), .C1(\U3/U12/DATA3_21 ), .C2(n870), .ZN(n100) );
  AOI22_X2 U301 ( .A1(\U3/U12/DATA1_22 ), .A2(n905), .B1(DiagonalY[22]), .B2(
        n903), .ZN(n101) );
  AOI222_X1 U302 ( .A1(\U3/U12/DATA2_22 ), .A2(n869), .B1(\U3/U12/DATA4_22 ), 
        .B2(n867), .C1(\U3/U12/DATA3_22 ), .C2(n870), .ZN(n102) );
  AOI22_X2 U304 ( .A1(\U3/U12/DATA1_23 ), .A2(n905), .B1(DiagonalY[23]), .B2(
        n903), .ZN(n103) );
  AOI222_X1 U305 ( .A1(\U3/U12/DATA2_23 ), .A2(n869), .B1(\U3/U12/DATA4_23 ), 
        .B2(n867), .C1(\U3/U12/DATA3_23 ), .C2(n870), .ZN(n104) );
  AOI22_X2 U307 ( .A1(\U3/U12/DATA1_24 ), .A2(n905), .B1(DiagonalY[24]), .B2(
        n903), .ZN(n105) );
  AOI222_X1 U308 ( .A1(\U3/U12/DATA2_24 ), .A2(n869), .B1(\U3/U12/DATA4_24 ), 
        .B2(n867), .C1(\U3/U12/DATA3_24 ), .C2(n870), .ZN(n106) );
  AOI22_X2 U310 ( .A1(\U3/U12/DATA1_25 ), .A2(n905), .B1(DiagonalY[25]), .B2(
        n903), .ZN(n107) );
  AOI222_X1 U311 ( .A1(\U3/U12/DATA2_25 ), .A2(n869), .B1(\U3/U12/DATA4_25 ), 
        .B2(n867), .C1(\U3/U12/DATA3_25 ), .C2(n870), .ZN(n108) );
  AOI22_X2 U313 ( .A1(\U3/U12/DATA1_26 ), .A2(n905), .B1(DiagonalY[26]), .B2(
        n903), .ZN(n109) );
  AOI222_X1 U314 ( .A1(\U3/U12/DATA2_26 ), .A2(n869), .B1(\U3/U12/DATA4_26 ), 
        .B2(n867), .C1(\U3/U12/DATA3_26 ), .C2(n870), .ZN(n110) );
  AOI22_X2 U316 ( .A1(\U3/U12/DATA1_27 ), .A2(n905), .B1(DiagonalY[27]), .B2(
        n903), .ZN(n111) );
  AOI222_X1 U317 ( .A1(\U3/U12/DATA2_27 ), .A2(n869), .B1(\U3/U12/DATA4_27 ), 
        .B2(n867), .C1(\U3/U12/DATA3_27 ), .C2(n870), .ZN(n112) );
  AOI22_X2 U319 ( .A1(\U3/U12/DATA1_28 ), .A2(n905), .B1(DiagonalY[28]), .B2(
        n903), .ZN(n113) );
  AOI222_X1 U320 ( .A1(\U3/U12/DATA2_28 ), .A2(n869), .B1(\U3/U12/DATA4_28 ), 
        .B2(n867), .C1(\U3/U12/DATA3_28 ), .C2(n870), .ZN(n114) );
  AOI22_X2 U322 ( .A1(\U3/U12/DATA1_29 ), .A2(n905), .B1(DiagonalY[29]), .B2(
        n903), .ZN(n115) );
  AOI222_X1 U323 ( .A1(\U3/U12/DATA2_29 ), .A2(n869), .B1(\U3/U12/DATA4_29 ), 
        .B2(n867), .C1(\U3/U12/DATA3_29 ), .C2(n870), .ZN(n116) );
  AOI22_X2 U325 ( .A1(\U3/U12/DATA1_30 ), .A2(n905), .B1(DiagonalY[30]), .B2(
        n903), .ZN(n117) );
  AOI222_X1 U326 ( .A1(\U3/U12/DATA2_30 ), .A2(n869), .B1(\U3/U12/DATA4_30 ), 
        .B2(n867), .C1(\U3/U12/DATA3_30 ), .C2(n870), .ZN(n118) );
  AOI22_X2 U328 ( .A1(\U3/U12/DATA1_31 ), .A2(n905), .B1(DiagonalY[31]), .B2(
        n903), .ZN(n119) );
  AOI222_X1 U329 ( .A1(\U3/U12/DATA2_31 ), .A2(n869), .B1(\U3/U12/DATA4_31 ), 
        .B2(n867), .C1(\U3/U12/DATA3_31 ), .C2(n870), .ZN(n120) );
  AOI22_X2 U331 ( .A1(\U3/U12/DATA1_32 ), .A2(n905), .B1(DiagonalY[32]), .B2(
        n903), .ZN(n121) );
  AOI222_X1 U332 ( .A1(\U3/U12/DATA2_32 ), .A2(n869), .B1(\U3/U12/DATA4_32 ), 
        .B2(n867), .C1(\U3/U12/DATA3_32 ), .C2(n870), .ZN(n122) );
  AOI22_X2 U334 ( .A1(\U3/U12/DATA1_33 ), .A2(n905), .B1(DiagonalY[33]), .B2(
        n903), .ZN(n123) );
  AOI222_X1 U335 ( .A1(\U3/U12/DATA2_33 ), .A2(n869), .B1(\U3/U12/DATA4_33 ), 
        .B2(n867), .C1(\U3/U12/DATA3_33 ), .C2(n870), .ZN(n124) );
  AOI22_X2 U337 ( .A1(\U3/U12/DATA1_34 ), .A2(n905), .B1(DiagonalY[34]), .B2(
        n903), .ZN(n125) );
  AOI222_X1 U338 ( .A1(\U3/U12/DATA2_34 ), .A2(n869), .B1(\U3/U12/DATA4_34 ), 
        .B2(n867), .C1(\U3/U12/DATA3_34 ), .C2(n870), .ZN(n126) );
  AOI22_X2 U340 ( .A1(\U3/U12/DATA1_35 ), .A2(n905), .B1(DiagonalY[35]), .B2(
        n903), .ZN(n127) );
  AOI222_X1 U341 ( .A1(\U3/U12/DATA2_35 ), .A2(n869), .B1(\U3/U12/DATA4_35 ), 
        .B2(n867), .C1(\U3/U12/DATA3_35 ), .C2(n870), .ZN(n128) );
  AOI22_X2 U343 ( .A1(\U3/U12/DATA1_36 ), .A2(n905), .B1(DiagonalY[36]), .B2(
        n903), .ZN(n129) );
  AOI222_X1 U344 ( .A1(\U3/U12/DATA2_36 ), .A2(n869), .B1(\U3/U12/DATA4_36 ), 
        .B2(n867), .C1(\U3/U12/DATA3_36 ), .C2(n870), .ZN(n130) );
  AOI22_X2 U346 ( .A1(\U3/U12/DATA1_37 ), .A2(n905), .B1(DiagonalY[37]), .B2(
        n903), .ZN(n131) );
  AOI222_X1 U347 ( .A1(\U3/U12/DATA2_37 ), .A2(n869), .B1(\U3/U12/DATA4_37 ), 
        .B2(n867), .C1(\U3/U12/DATA3_37 ), .C2(n870), .ZN(n132) );
  AOI22_X2 U349 ( .A1(\U3/U12/DATA1_38 ), .A2(n905), .B1(DiagonalY[38]), .B2(
        n903), .ZN(n133) );
  AOI222_X1 U350 ( .A1(\U3/U12/DATA2_38 ), .A2(n869), .B1(\U3/U12/DATA4_38 ), 
        .B2(n867), .C1(\U3/U12/DATA3_38 ), .C2(n870), .ZN(n134) );
  AOI22_X2 U352 ( .A1(\U3/U12/DATA1_39 ), .A2(n905), .B1(DiagonalY[39]), .B2(
        n903), .ZN(n135) );
  AOI222_X1 U353 ( .A1(\U3/U12/DATA2_39 ), .A2(n869), .B1(\U3/U12/DATA4_39 ), 
        .B2(n867), .C1(\U3/U12/DATA3_39 ), .C2(n870), .ZN(n136) );
  AOI22_X2 U355 ( .A1(\U3/U12/DATA1_40 ), .A2(n905), .B1(DiagonalY[40]), .B2(
        n903), .ZN(n137) );
  AOI222_X1 U356 ( .A1(\U3/U12/DATA2_40 ), .A2(n869), .B1(\U3/U12/DATA4_40 ), 
        .B2(n867), .C1(\U3/U12/DATA3_40 ), .C2(n870), .ZN(n138) );
  AOI22_X2 U358 ( .A1(\U3/U12/DATA1_41 ), .A2(n905), .B1(DiagonalY[41]), .B2(
        n903), .ZN(n139) );
  AOI222_X1 U359 ( .A1(\U3/U12/DATA2_41 ), .A2(n869), .B1(\U3/U12/DATA4_41 ), 
        .B2(n867), .C1(\U3/U12/DATA3_41 ), .C2(n870), .ZN(n140) );
  AOI22_X2 U361 ( .A1(\U3/U12/DATA1_42 ), .A2(n905), .B1(DiagonalY[42]), .B2(
        n903), .ZN(n141) );
  AOI222_X1 U362 ( .A1(\U3/U12/DATA2_42 ), .A2(n869), .B1(\U3/U12/DATA4_42 ), 
        .B2(n867), .C1(\U3/U12/DATA3_42 ), .C2(n870), .ZN(n142) );
  AOI22_X2 U364 ( .A1(\U3/U12/DATA1_43 ), .A2(n905), .B1(DiagonalY[43]), .B2(
        n903), .ZN(n143) );
  AOI222_X1 U365 ( .A1(\U3/U12/DATA2_43 ), .A2(n869), .B1(\U3/U12/DATA4_43 ), 
        .B2(n867), .C1(\U3/U12/DATA3_43 ), .C2(n870), .ZN(n144) );
  AOI22_X2 U367 ( .A1(\U3/U12/DATA1_44 ), .A2(n905), .B1(DiagonalY[44]), .B2(
        n903), .ZN(n145) );
  AOI222_X1 U368 ( .A1(\U3/U12/DATA2_44 ), .A2(n869), .B1(\U3/U12/DATA4_44 ), 
        .B2(n867), .C1(\U3/U12/DATA3_44 ), .C2(n870), .ZN(n146) );
  AOI22_X2 U370 ( .A1(\U3/U12/DATA1_45 ), .A2(n905), .B1(DiagonalY[45]), .B2(
        n903), .ZN(n147) );
  AOI222_X1 U371 ( .A1(\U3/U12/DATA2_45 ), .A2(n869), .B1(\U3/U12/DATA4_45 ), 
        .B2(n867), .C1(\U3/U12/DATA3_45 ), .C2(n870), .ZN(n148) );
  AOI22_X2 U373 ( .A1(\U3/U12/DATA1_46 ), .A2(n905), .B1(DiagonalY[46]), .B2(
        n903), .ZN(n149) );
  AOI222_X1 U374 ( .A1(\U3/U12/DATA2_46 ), .A2(n869), .B1(\U3/U12/DATA4_46 ), 
        .B2(n867), .C1(\U3/U12/DATA3_46 ), .C2(n870), .ZN(n150) );
  AOI22_X2 U376 ( .A1(\U3/U12/DATA1_47 ), .A2(n905), .B1(DiagonalY[47]), .B2(
        n903), .ZN(n151) );
  AOI222_X1 U377 ( .A1(\U3/U12/DATA2_47 ), .A2(n869), .B1(\U3/U12/DATA4_47 ), 
        .B2(n867), .C1(\U3/U12/DATA3_47 ), .C2(n870), .ZN(n152) );
  AOI22_X2 U379 ( .A1(PosDX[3]), .A2(n900), .B1(Row_noX[1]), .B2(n208), .ZN(
        n209) );
  AOI22_X2 U381 ( .A1(PosDX[4]), .A2(n900), .B1(Row_noX[2]), .B2(n208), .ZN(
        n210) );
  AOI22_X2 U382 ( .A1(PosDX[5]), .A2(n900), .B1(Row_noX[3]), .B2(n208), .ZN(
        n211) );
  AOI22_X2 U383 ( .A1(PosDX[6]), .A2(n900), .B1(Row_noX[4]), .B2(n208), .ZN(
        n212) );
  AOI22_X2 U436 ( .A1(PosDX[7]), .A2(n900), .B1(Row_noX[5]), .B2(n208), .ZN(
        n213) );
  AOI22_X2 U437 ( .A1(PosDX[8]), .A2(n900), .B1(Row_noX[6]), .B2(n208), .ZN(
        n214) );
  AOI22_X2 U438 ( .A1(PosDX[9]), .A2(n900), .B1(Row_noX[7]), .B2(n208), .ZN(
        n215) );
  AOI22_X2 U439 ( .A1(PosDX[10]), .A2(n900), .B1(Row_noX[8]), .B2(n208), .ZN(
        n216) );
  AOI22_X2 U440 ( .A1(PosDX[11]), .A2(n900), .B1(Row_noX[9]), .B2(n208), .ZN(
        n217) );
  AOI22_X2 U441 ( .A1(PosDX[2]), .A2(n900), .B1(Row_noX[0]), .B2(n208), .ZN(
        n207) );
  AOI22_X2 U442 ( .A1(PosDX[12]), .A2(n900), .B1(Row_noX[10]), .B2(n208), .ZN(
        n218) );
  INV_X4 U443 ( .A(n218), .ZN(n877) );
  INV_X4 U444 ( .A(n217), .ZN(n878) );
  INV_X4 U445 ( .A(n216), .ZN(n879) );
  INV_X4 U446 ( .A(n215), .ZN(n880) );
  INV_X4 U447 ( .A(n214), .ZN(n881) );
  INV_X4 U448 ( .A(n213), .ZN(n882) );
  INV_X4 U449 ( .A(n212), .ZN(n883) );
  INV_X4 U450 ( .A(n211), .ZN(n884) );
  INV_X4 U451 ( .A(n210), .ZN(n885) );
  INV_X4 U452 ( .A(n209), .ZN(n886) );
  INV_X4 U453 ( .A(n207), .ZN(n887) );
  INV_X4 U454 ( .A(n52), .ZN(n888) );
  INV_X4 U455 ( .A(n51), .ZN(n889) );
  INV_X4 U456 ( .A(n50), .ZN(n890) );
  INV_X4 U457 ( .A(n49), .ZN(n891) );
  INV_X4 U458 ( .A(n48), .ZN(n892) );
  INV_X4 U459 ( .A(n47), .ZN(n893) );
  INV_X4 U460 ( .A(n46), .ZN(n894) );
  INV_X4 U461 ( .A(n45), .ZN(n895) );
  INV_X4 U462 ( .A(n44), .ZN(n896) );
  INV_X4 U463 ( .A(n43), .ZN(n897) );
  INV_X4 U464 ( .A(n41), .ZN(n898) );
  INV_X4 U465 ( .A(n154), .ZN(n901) );
  INV_X4 U466 ( .A(n220), .ZN(n902) );
  INV_X4 U467 ( .A(n54), .ZN(n903) );
  INV_X4 U468 ( .A(n202), .ZN(n904) );
  INV_X4 U469 ( .A(n37), .ZN(n905) );
  INV_X4 U470 ( .A(n36), .ZN(n906) );
endmodule


module update_3_1 ( reset, clock, X, Y, NewRowX, NewRowY, Element, PosRowX, 
        PosRowY, PosDX, PosDY, FoundX, FoundY, Row_noX, Row_noY, DiagonalDoneX, 
        DiagonalDoneY, EnableChange, WireX, WireY );
  input [15:0] X;
  input [15:0] Y;
  input [255:0] NewRowX;
  input [255:0] NewRowY;
  output [47:0] Element;
  output [12:0] PosRowX;
  output [12:0] PosRowY;
  input [12:0] PosDX;
  input [12:0] PosDY;
  output [1:0] FoundX;
  output [1:0] FoundY;
  input [10:0] Row_noX;
  input [10:0] Row_noY;
  input reset, clock, DiagonalDoneX, DiagonalDoneY, EnableChange;
  output WireX, WireY;
  wire   \U168/DATA1_0 , \U168/DATA1_1 , \U168/DATA1_2 , \U168/DATA1_3 ,
         \U168/DATA1_4 , \U168/DATA1_5 , \U168/DATA1_6 , \U168/DATA1_7 ,
         \U168/DATA1_8 , \U168/DATA1_9 , \U168/DATA1_10 , \U168/DATA1_11 ,
         \U168/DATA1_12 , \U168/DATA1_13 , \U168/DATA1_14 , \U168/DATA1_15 ,
         \U168/DATA1_16 , \U168/DATA1_17 , \U168/DATA1_18 , \U168/DATA1_19 ,
         \U168/DATA1_20 , \U168/DATA1_21 , \U168/DATA1_22 , \U168/DATA1_23 ,
         \U168/DATA1_24 , \U168/DATA1_25 , \U168/DATA1_26 , \U168/DATA1_27 ,
         \U168/DATA1_28 , \U168/DATA1_29 , \U168/DATA1_30 , \U168/DATA1_31 ,
         \U168/DATA1_32 , \U168/DATA1_33 , \U168/DATA1_34 , \U168/DATA1_35 ,
         \U168/DATA1_36 , \U168/DATA1_37 , \U168/DATA1_38 , \U168/DATA1_39 ,
         \U168/DATA1_40 , \U168/DATA1_41 , \U168/DATA1_42 , \U168/DATA1_43 ,
         \U168/DATA1_44 , \U168/DATA1_45 , \U168/DATA1_46 , \U168/DATA1_47 ,
         \U166/DATA1_0 , \U166/DATA1_1 , \U166/DATA1_2 , \U166/DATA1_3 ,
         \U166/DATA1_4 , \U166/DATA1_5 , \U166/DATA1_6 , \U166/DATA1_7 ,
         \U166/DATA1_8 , \U166/DATA1_9 , \U166/DATA1_10 , \U166/DATA1_11 ,
         \U166/DATA1_12 , \U166/DATA1_13 , \U166/DATA1_14 , \U166/DATA1_15 ,
         \U166/DATA1_16 , \U166/DATA1_17 , \U166/DATA1_18 , \U166/DATA1_19 ,
         \U166/DATA1_20 , \U166/DATA1_21 , \U166/DATA1_22 , \U166/DATA1_23 ,
         \U166/DATA1_24 , \U166/DATA1_25 , \U166/DATA1_26 , \U166/DATA1_27 ,
         \U166/DATA1_28 , \U166/DATA1_29 , \U166/DATA1_30 , \U166/DATA1_31 ,
         \U166/DATA1_32 , \U166/DATA1_33 , \U166/DATA1_34 , \U166/DATA1_35 ,
         \U166/DATA1_36 , \U166/DATA1_37 , \U166/DATA1_38 , \U166/DATA1_39 ,
         \U166/DATA1_40 , \U166/DATA1_41 , \U166/DATA1_42 , \U166/DATA1_43 ,
         \U166/DATA1_44 , \U166/DATA1_45 , \U166/DATA1_46 , \U166/DATA1_47 ,
         \U163/DATA1_0 , \U163/DATA1_1 , \U163/DATA1_2 , \U163/DATA1_3 ,
         \U163/DATA1_4 , \U163/DATA1_5 , \U163/DATA1_6 , \U163/DATA1_7 ,
         \U163/DATA1_8 , \U163/DATA1_9 , \U163/DATA1_10 , \U163/DATA1_11 ,
         \U163/DATA1_12 , \U163/DATA1_13 , \U163/DATA1_14 , \U163/DATA1_15 ,
         \U163/DATA1_16 , \U163/DATA1_17 , \U163/DATA1_18 , \U163/DATA1_19 ,
         \U163/DATA1_20 , \U163/DATA1_21 , \U163/DATA1_22 , \U163/DATA1_23 ,
         \U163/DATA1_24 , \U163/DATA1_25 , \U163/DATA1_26 , \U163/DATA1_27 ,
         \U163/DATA1_28 , \U163/DATA1_29 , \U163/DATA1_30 , \U163/DATA1_31 ,
         \U163/DATA1_32 , \U163/DATA1_33 , \U163/DATA1_34 , \U163/DATA1_35 ,
         \U163/DATA1_36 , \U163/DATA1_37 , \U163/DATA1_38 , \U163/DATA1_39 ,
         \U163/DATA1_40 , \U163/DATA1_41 , \U163/DATA1_42 , \U163/DATA1_43 ,
         \U163/DATA1_44 , \U163/DATA1_45 , \U163/DATA1_46 , \U163/DATA1_47 ,
         \U125/DATA1_0 , \U125/DATA1_1 , \U125/DATA1_2 , \U125/DATA1_3 ,
         \U125/DATA1_4 , \U125/DATA1_5 , \U125/DATA1_6 , \U125/DATA1_7 ,
         \U125/DATA1_8 , \U125/DATA1_9 , \U125/DATA1_10 , \U125/DATA1_11 ,
         \U125/DATA1_12 , \U125/DATA1_13 , \U125/DATA1_14 , \U125/DATA1_15 ,
         \U125/DATA1_16 , \U125/DATA1_17 , \U125/DATA1_18 , \U125/DATA1_19 ,
         \U125/DATA1_20 , \U125/DATA1_21 , \U125/DATA1_22 , \U125/DATA1_23 ,
         \U125/DATA1_24 , \U125/DATA1_25 , \U125/DATA1_26 , \U125/DATA1_27 ,
         \U125/DATA1_28 , \U125/DATA1_29 , \U125/DATA1_30 , \U125/DATA1_31 ,
         \U125/DATA1_32 , \U125/DATA1_33 , \U125/DATA1_34 , \U125/DATA1_35 ,
         \U125/DATA1_36 , \U125/DATA1_37 , \U125/DATA1_38 , \U125/DATA1_39 ,
         \U125/DATA1_40 , \U125/DATA1_41 , \U125/DATA1_42 , \U125/DATA1_43 ,
         \U125/DATA1_44 , \U125/DATA1_45 , \U125/DATA1_46 , \U125/DATA1_47 ,
         \U95/DATA1_0 , \U95/DATA1_1 , \U95/DATA1_2 , \U95/DATA1_3 ,
         \U95/DATA1_4 , \U95/DATA1_5 , \U95/DATA1_6 , \U95/DATA1_7 ,
         \U95/DATA1_8 , \U95/DATA1_9 , \U95/DATA1_10 , \U95/DATA1_11 ,
         \U95/DATA1_12 , \U95/DATA1_13 , \U95/DATA1_14 , \U95/DATA1_15 ,
         \U95/DATA1_16 , \U95/DATA1_17 , \U95/DATA1_18 , \U95/DATA1_19 ,
         \U95/DATA1_20 , \U95/DATA1_21 , \U95/DATA1_22 , \U95/DATA1_23 ,
         \U95/DATA1_24 , \U95/DATA1_25 , \U95/DATA1_26 , \U95/DATA1_27 ,
         \U95/DATA1_28 , \U95/DATA1_29 , \U95/DATA1_30 , \U95/DATA1_31 ,
         \U95/DATA1_32 , \U95/DATA1_33 , \U95/DATA1_34 , \U95/DATA1_35 ,
         \U95/DATA1_36 , \U95/DATA1_37 , \U95/DATA1_38 , \U95/DATA1_39 ,
         \U95/DATA1_40 , \U95/DATA1_41 , \U95/DATA1_42 , \U95/DATA1_43 ,
         \U95/DATA1_44 , \U95/DATA1_45 , \U95/DATA1_46 , \U95/DATA1_47 ,
         \U93/DATA1_0 , \U93/DATA1_1 , \U93/DATA1_2 , \U93/DATA1_3 ,
         \U93/DATA1_4 , \U93/DATA1_5 , \U93/DATA1_6 , \U93/DATA1_7 ,
         \U93/DATA1_8 , \U93/DATA1_9 , \U93/DATA1_10 , \U93/DATA1_11 ,
         \U93/DATA1_12 , \U93/DATA1_13 , \U93/DATA1_14 , \U93/DATA1_15 ,
         \U93/DATA1_16 , \U93/DATA1_17 , \U93/DATA1_18 , \U93/DATA1_19 ,
         \U93/DATA1_20 , \U93/DATA1_21 , \U93/DATA1_22 , \U93/DATA1_23 ,
         \U93/DATA1_24 , \U93/DATA1_25 , \U93/DATA1_26 , \U93/DATA1_27 ,
         \U93/DATA1_28 , \U93/DATA1_29 , \U93/DATA1_30 , \U93/DATA1_31 ,
         \U93/DATA1_32 , \U93/DATA1_33 , \U93/DATA1_34 , \U93/DATA1_35 ,
         \U93/DATA1_36 , \U93/DATA1_37 , \U93/DATA1_38 , \U93/DATA1_39 ,
         \U93/DATA1_40 , \U93/DATA1_41 , \U93/DATA1_42 , \U93/DATA1_43 ,
         \U93/DATA1_44 , \U93/DATA1_45 , \U93/DATA1_46 , \U93/DATA1_47 ,
         \U90/DATA1_0 , \U90/DATA1_1 , \U90/DATA1_2 , \U90/DATA1_3 ,
         \U90/DATA1_4 , \U90/DATA1_5 , \U90/DATA1_6 , \U90/DATA1_7 ,
         \U90/DATA1_8 , \U90/DATA1_9 , \U90/DATA1_10 , \U90/DATA1_11 ,
         \U90/DATA1_12 , \U90/DATA1_13 , \U90/DATA1_14 , \U90/DATA1_15 ,
         \U90/DATA1_16 , \U90/DATA1_17 , \U90/DATA1_18 , \U90/DATA1_19 ,
         \U90/DATA1_20 , \U90/DATA1_21 , \U90/DATA1_22 , \U90/DATA1_23 ,
         \U90/DATA1_24 , \U90/DATA1_25 , \U90/DATA1_26 , \U90/DATA1_27 ,
         \U90/DATA1_28 , \U90/DATA1_29 , \U90/DATA1_30 , \U90/DATA1_31 ,
         \U90/DATA1_32 , \U90/DATA1_33 , \U90/DATA1_34 , \U90/DATA1_35 ,
         \U90/DATA1_36 , \U90/DATA1_37 , \U90/DATA1_38 , \U90/DATA1_39 ,
         \U90/DATA1_40 , \U90/DATA1_41 , \U90/DATA1_42 , \U90/DATA1_43 ,
         \U90/DATA1_44 , \U90/DATA1_45 , \U90/DATA1_46 , \U90/DATA1_47 ,
         \U52/DATA1_0 , \U52/DATA1_1 , \U52/DATA1_2 , \U52/DATA1_3 ,
         \U52/DATA1_4 , \U52/DATA1_5 , \U52/DATA1_6 , \U52/DATA1_7 ,
         \U52/DATA1_8 , \U52/DATA1_9 , \U52/DATA1_10 , \U52/DATA1_11 ,
         \U52/DATA1_12 , \U52/DATA1_13 , \U52/DATA1_14 , \U52/DATA1_15 ,
         \U52/DATA1_16 , \U52/DATA1_17 , \U52/DATA1_18 , \U52/DATA1_19 ,
         \U52/DATA1_20 , \U52/DATA1_21 , \U52/DATA1_22 , \U52/DATA1_23 ,
         \U52/DATA1_24 , \U52/DATA1_25 , \U52/DATA1_26 , \U52/DATA1_27 ,
         \U52/DATA1_28 , \U52/DATA1_29 , \U52/DATA1_30 , \U52/DATA1_31 ,
         \U52/DATA1_32 , \U52/DATA1_33 , \U52/DATA1_34 , \U52/DATA1_35 ,
         \U52/DATA1_36 , \U52/DATA1_37 , \U52/DATA1_38 , \U52/DATA1_39 ,
         \U52/DATA1_40 , \U52/DATA1_41 , \U52/DATA1_42 , \U52/DATA1_43 ,
         \U52/DATA1_44 , \U52/DATA1_45 , \U52/DATA1_46 , \U52/DATA1_47 ,
         \eq_207/A[15] , \eq_207/A[14] , \eq_207/A[13] , \eq_207/A[12] ,
         \eq_207/A[11] , \eq_207/A[10] , \eq_207/A[9] , \eq_207/A[8] ,
         \eq_207/A[7] , \eq_207/A[6] , \eq_207/A[5] , \eq_207/A[4] ,
         \eq_207/A[3] , \eq_207/A[2] , \eq_207/A[1] , \eq_207/A[0] ,
         \eq_207/B[15] , \eq_207/B[14] , \eq_207/B[13] , \eq_207/B[12] ,
         \eq_207/B[11] , \eq_207/B[10] , \eq_207/B[9] , \eq_207/B[8] ,
         \eq_207/B[7] , \eq_207/B[6] , \eq_207/B[5] , \eq_207/B[4] ,
         \eq_207/B[3] , \eq_207/B[2] , \eq_207/B[1] , \eq_207/B[0] ,
         \eq_112/A[15] , \eq_112/A[14] , \eq_112/A[13] , \eq_112/A[12] ,
         \eq_112/A[11] , \eq_112/A[10] , \eq_112/A[9] , \eq_112/A[8] ,
         \eq_112/A[7] , \eq_112/A[6] , \eq_112/A[5] , \eq_112/A[4] ,
         \eq_112/A[3] , \eq_112/A[2] , \eq_112/A[1] , \eq_112/A[0] ,
         \eq_112/B[15] , \eq_112/B[14] , \eq_112/B[13] , \eq_112/B[12] ,
         \eq_112/B[11] , \eq_112/B[10] , \eq_112/B[9] , \eq_112/B[8] ,
         \eq_112/B[7] , \eq_112/B[6] , \eq_112/B[5] , \eq_112/B[4] ,
         \eq_112/B[3] , \eq_112/B[2] , \eq_112/B[1] , \eq_112/B[0] ,
         \r528/A[15] , \r528/A[14] , \r528/A[13] , \r528/A[12] , \r528/A[11] ,
         \r528/A[10] , \r528/A[9] , \r528/A[8] , \r528/A[7] , \r528/A[6] ,
         \r528/A[5] , \r528/A[4] , \r528/A[3] , \r528/A[2] , \r528/A[1] ,
         \r528/A[0] , \r527/A[15] , \r527/A[14] , \r527/A[13] , \r527/A[12] ,
         \r527/A[11] , \r527/A[10] , \r527/A[9] , \r527/A[8] , \r527/A[7] ,
         \r527/A[6] , \r527/A[5] , \r527/A[4] , \r527/A[3] , \r527/A[2] ,
         \r527/A[1] , \r527/A[0] , \r526/A[15] , \r526/A[14] , \r526/A[13] ,
         \r526/A[12] , \r526/A[11] , \r526/A[10] , \r526/A[9] , \r526/A[8] ,
         \r526/A[7] , \r526/A[6] , \r526/A[5] , \r526/A[4] , \r526/A[3] ,
         \r526/A[2] , \r526/A[1] , \r526/A[0] , \r524/A[15] , \r524/A[14] ,
         \r524/A[13] , \r524/A[12] , \r524/A[11] , \r524/A[10] , \r524/A[9] ,
         \r524/A[8] , \r524/A[7] , \r524/A[6] , \r524/A[5] , \r524/A[4] ,
         \r524/A[3] , \r524/A[2] , \r524/A[1] , \r524/A[0] , \r523/A[15] ,
         \r523/A[14] , \r523/A[13] , \r523/A[12] , \r523/A[11] , \r523/A[10] ,
         \r523/A[9] , \r523/A[8] , \r523/A[7] , \r523/A[6] , \r523/A[5] ,
         \r523/A[4] , \r523/A[3] , \r523/A[2] , \r523/A[1] , \r523/A[0] ,
         \r522/A[15] , \r522/A[14] , \r522/A[13] , \r522/A[12] , \r522/A[11] ,
         \r522/A[10] , \r522/A[9] , \r522/A[8] , \r522/A[7] , \r522/A[6] ,
         \r522/A[5] , \r522/A[4] , \r522/A[3] , \r522/A[2] , \r522/A[1] ,
         \r522/A[0] , n28, n29, n35, n36, n193, n194, n196, n197, n198, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n217, n218, n220, n221, n222, n223, n226,
         n228, n231, n232, n234, n235, n239, n242, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110;
  assign \U168/DATA1_0  = NewRowX[128];
  assign \U168/DATA1_1  = NewRowX[129];
  assign \U168/DATA1_2  = NewRowX[130];
  assign \U168/DATA1_3  = NewRowX[131];
  assign \U168/DATA1_4  = NewRowX[132];
  assign \U168/DATA1_5  = NewRowX[133];
  assign \U168/DATA1_6  = NewRowX[134];
  assign \U168/DATA1_7  = NewRowX[135];
  assign \U168/DATA1_8  = NewRowX[136];
  assign \U168/DATA1_9  = NewRowX[137];
  assign \U168/DATA1_10  = NewRowX[138];
  assign \U168/DATA1_11  = NewRowX[139];
  assign \U168/DATA1_12  = NewRowX[140];
  assign \U168/DATA1_13  = NewRowX[141];
  assign \U168/DATA1_14  = NewRowX[142];
  assign \U168/DATA1_15  = NewRowX[143];
  assign \U168/DATA1_16  = NewRowX[144];
  assign \U168/DATA1_17  = NewRowX[145];
  assign \U168/DATA1_18  = NewRowX[146];
  assign \U168/DATA1_19  = NewRowX[147];
  assign \U168/DATA1_20  = NewRowX[148];
  assign \U168/DATA1_21  = NewRowX[149];
  assign \U168/DATA1_22  = NewRowX[150];
  assign \U168/DATA1_23  = NewRowX[151];
  assign \U168/DATA1_24  = NewRowX[152];
  assign \U168/DATA1_25  = NewRowX[153];
  assign \U168/DATA1_26  = NewRowX[154];
  assign \U168/DATA1_27  = NewRowX[155];
  assign \U168/DATA1_28  = NewRowX[156];
  assign \U168/DATA1_29  = NewRowX[157];
  assign \U168/DATA1_30  = NewRowX[158];
  assign \U168/DATA1_31  = NewRowX[159];
  assign \U168/DATA1_32  = NewRowX[160];
  assign \U168/DATA1_33  = NewRowX[161];
  assign \U168/DATA1_34  = NewRowX[162];
  assign \U168/DATA1_35  = NewRowX[163];
  assign \U168/DATA1_36  = NewRowX[164];
  assign \U168/DATA1_37  = NewRowX[165];
  assign \U168/DATA1_38  = NewRowX[166];
  assign \U168/DATA1_39  = NewRowX[167];
  assign \U168/DATA1_40  = NewRowX[168];
  assign \U168/DATA1_41  = NewRowX[169];
  assign \U168/DATA1_42  = NewRowX[170];
  assign \U168/DATA1_43  = NewRowX[171];
  assign \U168/DATA1_44  = NewRowX[172];
  assign \U168/DATA1_45  = NewRowX[173];
  assign \U168/DATA1_46  = NewRowX[174];
  assign \U168/DATA1_47  = NewRowX[175];
  assign \U166/DATA1_0  = NewRowX[64];
  assign \U166/DATA1_1  = NewRowX[65];
  assign \U166/DATA1_2  = NewRowX[66];
  assign \U166/DATA1_3  = NewRowX[67];
  assign \U166/DATA1_4  = NewRowX[68];
  assign \U166/DATA1_5  = NewRowX[69];
  assign \U166/DATA1_6  = NewRowX[70];
  assign \U166/DATA1_7  = NewRowX[71];
  assign \U166/DATA1_8  = NewRowX[72];
  assign \U166/DATA1_9  = NewRowX[73];
  assign \U166/DATA1_10  = NewRowX[74];
  assign \U166/DATA1_11  = NewRowX[75];
  assign \U166/DATA1_12  = NewRowX[76];
  assign \U166/DATA1_13  = NewRowX[77];
  assign \U166/DATA1_14  = NewRowX[78];
  assign \U166/DATA1_15  = NewRowX[79];
  assign \U166/DATA1_16  = NewRowX[80];
  assign \U166/DATA1_17  = NewRowX[81];
  assign \U166/DATA1_18  = NewRowX[82];
  assign \U166/DATA1_19  = NewRowX[83];
  assign \U166/DATA1_20  = NewRowX[84];
  assign \U166/DATA1_21  = NewRowX[85];
  assign \U166/DATA1_22  = NewRowX[86];
  assign \U166/DATA1_23  = NewRowX[87];
  assign \U166/DATA1_24  = NewRowX[88];
  assign \U166/DATA1_25  = NewRowX[89];
  assign \U166/DATA1_26  = NewRowX[90];
  assign \U166/DATA1_27  = NewRowX[91];
  assign \U166/DATA1_28  = NewRowX[92];
  assign \U166/DATA1_29  = NewRowX[93];
  assign \U166/DATA1_30  = NewRowX[94];
  assign \U166/DATA1_31  = NewRowX[95];
  assign \U166/DATA1_32  = NewRowX[96];
  assign \U166/DATA1_33  = NewRowX[97];
  assign \U166/DATA1_34  = NewRowX[98];
  assign \U166/DATA1_35  = NewRowX[99];
  assign \U166/DATA1_36  = NewRowX[100];
  assign \U166/DATA1_37  = NewRowX[101];
  assign \U166/DATA1_38  = NewRowX[102];
  assign \U166/DATA1_39  = NewRowX[103];
  assign \U166/DATA1_40  = NewRowX[104];
  assign \U166/DATA1_41  = NewRowX[105];
  assign \U166/DATA1_42  = NewRowX[106];
  assign \U166/DATA1_43  = NewRowX[107];
  assign \U166/DATA1_44  = NewRowX[108];
  assign \U166/DATA1_45  = NewRowX[109];
  assign \U166/DATA1_46  = NewRowX[110];
  assign \U166/DATA1_47  = NewRowX[111];
  assign \U163/DATA1_0  = NewRowX[0];
  assign \U163/DATA1_1  = NewRowX[1];
  assign \U163/DATA1_2  = NewRowX[2];
  assign \U163/DATA1_3  = NewRowX[3];
  assign \U163/DATA1_4  = NewRowX[4];
  assign \U163/DATA1_5  = NewRowX[5];
  assign \U163/DATA1_6  = NewRowX[6];
  assign \U163/DATA1_7  = NewRowX[7];
  assign \U163/DATA1_8  = NewRowX[8];
  assign \U163/DATA1_9  = NewRowX[9];
  assign \U163/DATA1_10  = NewRowX[10];
  assign \U163/DATA1_11  = NewRowX[11];
  assign \U163/DATA1_12  = NewRowX[12];
  assign \U163/DATA1_13  = NewRowX[13];
  assign \U163/DATA1_14  = NewRowX[14];
  assign \U163/DATA1_15  = NewRowX[15];
  assign \U163/DATA1_16  = NewRowX[16];
  assign \U163/DATA1_17  = NewRowX[17];
  assign \U163/DATA1_18  = NewRowX[18];
  assign \U163/DATA1_19  = NewRowX[19];
  assign \U163/DATA1_20  = NewRowX[20];
  assign \U163/DATA1_21  = NewRowX[21];
  assign \U163/DATA1_22  = NewRowX[22];
  assign \U163/DATA1_23  = NewRowX[23];
  assign \U163/DATA1_24  = NewRowX[24];
  assign \U163/DATA1_25  = NewRowX[25];
  assign \U163/DATA1_26  = NewRowX[26];
  assign \U163/DATA1_27  = NewRowX[27];
  assign \U163/DATA1_28  = NewRowX[28];
  assign \U163/DATA1_29  = NewRowX[29];
  assign \U163/DATA1_30  = NewRowX[30];
  assign \U163/DATA1_31  = NewRowX[31];
  assign \U163/DATA1_32  = NewRowX[32];
  assign \U163/DATA1_33  = NewRowX[33];
  assign \U163/DATA1_34  = NewRowX[34];
  assign \U163/DATA1_35  = NewRowX[35];
  assign \U163/DATA1_36  = NewRowX[36];
  assign \U163/DATA1_37  = NewRowX[37];
  assign \U163/DATA1_38  = NewRowX[38];
  assign \U163/DATA1_39  = NewRowX[39];
  assign \U163/DATA1_40  = NewRowX[40];
  assign \U163/DATA1_41  = NewRowX[41];
  assign \U163/DATA1_42  = NewRowX[42];
  assign \U163/DATA1_43  = NewRowX[43];
  assign \U163/DATA1_44  = NewRowX[44];
  assign \U163/DATA1_45  = NewRowX[45];
  assign \U163/DATA1_46  = NewRowX[46];
  assign \U163/DATA1_47  = NewRowX[47];
  assign \U125/DATA1_0  = NewRowX[192];
  assign \U125/DATA1_1  = NewRowX[193];
  assign \U125/DATA1_2  = NewRowX[194];
  assign \U125/DATA1_3  = NewRowX[195];
  assign \U125/DATA1_4  = NewRowX[196];
  assign \U125/DATA1_5  = NewRowX[197];
  assign \U125/DATA1_6  = NewRowX[198];
  assign \U125/DATA1_7  = NewRowX[199];
  assign \U125/DATA1_8  = NewRowX[200];
  assign \U125/DATA1_9  = NewRowX[201];
  assign \U125/DATA1_10  = NewRowX[202];
  assign \U125/DATA1_11  = NewRowX[203];
  assign \U125/DATA1_12  = NewRowX[204];
  assign \U125/DATA1_13  = NewRowX[205];
  assign \U125/DATA1_14  = NewRowX[206];
  assign \U125/DATA1_15  = NewRowX[207];
  assign \U125/DATA1_16  = NewRowX[208];
  assign \U125/DATA1_17  = NewRowX[209];
  assign \U125/DATA1_18  = NewRowX[210];
  assign \U125/DATA1_19  = NewRowX[211];
  assign \U125/DATA1_20  = NewRowX[212];
  assign \U125/DATA1_21  = NewRowX[213];
  assign \U125/DATA1_22  = NewRowX[214];
  assign \U125/DATA1_23  = NewRowX[215];
  assign \U125/DATA1_24  = NewRowX[216];
  assign \U125/DATA1_25  = NewRowX[217];
  assign \U125/DATA1_26  = NewRowX[218];
  assign \U125/DATA1_27  = NewRowX[219];
  assign \U125/DATA1_28  = NewRowX[220];
  assign \U125/DATA1_29  = NewRowX[221];
  assign \U125/DATA1_30  = NewRowX[222];
  assign \U125/DATA1_31  = NewRowX[223];
  assign \U125/DATA1_32  = NewRowX[224];
  assign \U125/DATA1_33  = NewRowX[225];
  assign \U125/DATA1_34  = NewRowX[226];
  assign \U125/DATA1_35  = NewRowX[227];
  assign \U125/DATA1_36  = NewRowX[228];
  assign \U125/DATA1_37  = NewRowX[229];
  assign \U125/DATA1_38  = NewRowX[230];
  assign \U125/DATA1_39  = NewRowX[231];
  assign \U125/DATA1_40  = NewRowX[232];
  assign \U125/DATA1_41  = NewRowX[233];
  assign \U125/DATA1_42  = NewRowX[234];
  assign \U125/DATA1_43  = NewRowX[235];
  assign \U125/DATA1_44  = NewRowX[236];
  assign \U125/DATA1_45  = NewRowX[237];
  assign \U125/DATA1_46  = NewRowX[238];
  assign \U125/DATA1_47  = NewRowX[239];
  assign \U95/DATA1_0  = NewRowY[128];
  assign \U95/DATA1_1  = NewRowY[129];
  assign \U95/DATA1_2  = NewRowY[130];
  assign \U95/DATA1_3  = NewRowY[131];
  assign \U95/DATA1_4  = NewRowY[132];
  assign \U95/DATA1_5  = NewRowY[133];
  assign \U95/DATA1_6  = NewRowY[134];
  assign \U95/DATA1_7  = NewRowY[135];
  assign \U95/DATA1_8  = NewRowY[136];
  assign \U95/DATA1_9  = NewRowY[137];
  assign \U95/DATA1_10  = NewRowY[138];
  assign \U95/DATA1_11  = NewRowY[139];
  assign \U95/DATA1_12  = NewRowY[140];
  assign \U95/DATA1_13  = NewRowY[141];
  assign \U95/DATA1_14  = NewRowY[142];
  assign \U95/DATA1_15  = NewRowY[143];
  assign \U95/DATA1_16  = NewRowY[144];
  assign \U95/DATA1_17  = NewRowY[145];
  assign \U95/DATA1_18  = NewRowY[146];
  assign \U95/DATA1_19  = NewRowY[147];
  assign \U95/DATA1_20  = NewRowY[148];
  assign \U95/DATA1_21  = NewRowY[149];
  assign \U95/DATA1_22  = NewRowY[150];
  assign \U95/DATA1_23  = NewRowY[151];
  assign \U95/DATA1_24  = NewRowY[152];
  assign \U95/DATA1_25  = NewRowY[153];
  assign \U95/DATA1_26  = NewRowY[154];
  assign \U95/DATA1_27  = NewRowY[155];
  assign \U95/DATA1_28  = NewRowY[156];
  assign \U95/DATA1_29  = NewRowY[157];
  assign \U95/DATA1_30  = NewRowY[158];
  assign \U95/DATA1_31  = NewRowY[159];
  assign \U95/DATA1_32  = NewRowY[160];
  assign \U95/DATA1_33  = NewRowY[161];
  assign \U95/DATA1_34  = NewRowY[162];
  assign \U95/DATA1_35  = NewRowY[163];
  assign \U95/DATA1_36  = NewRowY[164];
  assign \U95/DATA1_37  = NewRowY[165];
  assign \U95/DATA1_38  = NewRowY[166];
  assign \U95/DATA1_39  = NewRowY[167];
  assign \U95/DATA1_40  = NewRowY[168];
  assign \U95/DATA1_41  = NewRowY[169];
  assign \U95/DATA1_42  = NewRowY[170];
  assign \U95/DATA1_43  = NewRowY[171];
  assign \U95/DATA1_44  = NewRowY[172];
  assign \U95/DATA1_45  = NewRowY[173];
  assign \U95/DATA1_46  = NewRowY[174];
  assign \U95/DATA1_47  = NewRowY[175];
  assign \U93/DATA1_0  = NewRowY[64];
  assign \U93/DATA1_1  = NewRowY[65];
  assign \U93/DATA1_2  = NewRowY[66];
  assign \U93/DATA1_3  = NewRowY[67];
  assign \U93/DATA1_4  = NewRowY[68];
  assign \U93/DATA1_5  = NewRowY[69];
  assign \U93/DATA1_6  = NewRowY[70];
  assign \U93/DATA1_7  = NewRowY[71];
  assign \U93/DATA1_8  = NewRowY[72];
  assign \U93/DATA1_9  = NewRowY[73];
  assign \U93/DATA1_10  = NewRowY[74];
  assign \U93/DATA1_11  = NewRowY[75];
  assign \U93/DATA1_12  = NewRowY[76];
  assign \U93/DATA1_13  = NewRowY[77];
  assign \U93/DATA1_14  = NewRowY[78];
  assign \U93/DATA1_15  = NewRowY[79];
  assign \U93/DATA1_16  = NewRowY[80];
  assign \U93/DATA1_17  = NewRowY[81];
  assign \U93/DATA1_18  = NewRowY[82];
  assign \U93/DATA1_19  = NewRowY[83];
  assign \U93/DATA1_20  = NewRowY[84];
  assign \U93/DATA1_21  = NewRowY[85];
  assign \U93/DATA1_22  = NewRowY[86];
  assign \U93/DATA1_23  = NewRowY[87];
  assign \U93/DATA1_24  = NewRowY[88];
  assign \U93/DATA1_25  = NewRowY[89];
  assign \U93/DATA1_26  = NewRowY[90];
  assign \U93/DATA1_27  = NewRowY[91];
  assign \U93/DATA1_28  = NewRowY[92];
  assign \U93/DATA1_29  = NewRowY[93];
  assign \U93/DATA1_30  = NewRowY[94];
  assign \U93/DATA1_31  = NewRowY[95];
  assign \U93/DATA1_32  = NewRowY[96];
  assign \U93/DATA1_33  = NewRowY[97];
  assign \U93/DATA1_34  = NewRowY[98];
  assign \U93/DATA1_35  = NewRowY[99];
  assign \U93/DATA1_36  = NewRowY[100];
  assign \U93/DATA1_37  = NewRowY[101];
  assign \U93/DATA1_38  = NewRowY[102];
  assign \U93/DATA1_39  = NewRowY[103];
  assign \U93/DATA1_40  = NewRowY[104];
  assign \U93/DATA1_41  = NewRowY[105];
  assign \U93/DATA1_42  = NewRowY[106];
  assign \U93/DATA1_43  = NewRowY[107];
  assign \U93/DATA1_44  = NewRowY[108];
  assign \U93/DATA1_45  = NewRowY[109];
  assign \U93/DATA1_46  = NewRowY[110];
  assign \U93/DATA1_47  = NewRowY[111];
  assign \U90/DATA1_0  = NewRowY[0];
  assign \U90/DATA1_1  = NewRowY[1];
  assign \U90/DATA1_2  = NewRowY[2];
  assign \U90/DATA1_3  = NewRowY[3];
  assign \U90/DATA1_4  = NewRowY[4];
  assign \U90/DATA1_5  = NewRowY[5];
  assign \U90/DATA1_6  = NewRowY[6];
  assign \U90/DATA1_7  = NewRowY[7];
  assign \U90/DATA1_8  = NewRowY[8];
  assign \U90/DATA1_9  = NewRowY[9];
  assign \U90/DATA1_10  = NewRowY[10];
  assign \U90/DATA1_11  = NewRowY[11];
  assign \U90/DATA1_12  = NewRowY[12];
  assign \U90/DATA1_13  = NewRowY[13];
  assign \U90/DATA1_14  = NewRowY[14];
  assign \U90/DATA1_15  = NewRowY[15];
  assign \U90/DATA1_16  = NewRowY[16];
  assign \U90/DATA1_17  = NewRowY[17];
  assign \U90/DATA1_18  = NewRowY[18];
  assign \U90/DATA1_19  = NewRowY[19];
  assign \U90/DATA1_20  = NewRowY[20];
  assign \U90/DATA1_21  = NewRowY[21];
  assign \U90/DATA1_22  = NewRowY[22];
  assign \U90/DATA1_23  = NewRowY[23];
  assign \U90/DATA1_24  = NewRowY[24];
  assign \U90/DATA1_25  = NewRowY[25];
  assign \U90/DATA1_26  = NewRowY[26];
  assign \U90/DATA1_27  = NewRowY[27];
  assign \U90/DATA1_28  = NewRowY[28];
  assign \U90/DATA1_29  = NewRowY[29];
  assign \U90/DATA1_30  = NewRowY[30];
  assign \U90/DATA1_31  = NewRowY[31];
  assign \U90/DATA1_32  = NewRowY[32];
  assign \U90/DATA1_33  = NewRowY[33];
  assign \U90/DATA1_34  = NewRowY[34];
  assign \U90/DATA1_35  = NewRowY[35];
  assign \U90/DATA1_36  = NewRowY[36];
  assign \U90/DATA1_37  = NewRowY[37];
  assign \U90/DATA1_38  = NewRowY[38];
  assign \U90/DATA1_39  = NewRowY[39];
  assign \U90/DATA1_40  = NewRowY[40];
  assign \U90/DATA1_41  = NewRowY[41];
  assign \U90/DATA1_42  = NewRowY[42];
  assign \U90/DATA1_43  = NewRowY[43];
  assign \U90/DATA1_44  = NewRowY[44];
  assign \U90/DATA1_45  = NewRowY[45];
  assign \U90/DATA1_46  = NewRowY[46];
  assign \U90/DATA1_47  = NewRowY[47];
  assign \U52/DATA1_0  = NewRowY[192];
  assign \U52/DATA1_1  = NewRowY[193];
  assign \U52/DATA1_2  = NewRowY[194];
  assign \U52/DATA1_3  = NewRowY[195];
  assign \U52/DATA1_4  = NewRowY[196];
  assign \U52/DATA1_5  = NewRowY[197];
  assign \U52/DATA1_6  = NewRowY[198];
  assign \U52/DATA1_7  = NewRowY[199];
  assign \U52/DATA1_8  = NewRowY[200];
  assign \U52/DATA1_9  = NewRowY[201];
  assign \U52/DATA1_10  = NewRowY[202];
  assign \U52/DATA1_11  = NewRowY[203];
  assign \U52/DATA1_12  = NewRowY[204];
  assign \U52/DATA1_13  = NewRowY[205];
  assign \U52/DATA1_14  = NewRowY[206];
  assign \U52/DATA1_15  = NewRowY[207];
  assign \U52/DATA1_16  = NewRowY[208];
  assign \U52/DATA1_17  = NewRowY[209];
  assign \U52/DATA1_18  = NewRowY[210];
  assign \U52/DATA1_19  = NewRowY[211];
  assign \U52/DATA1_20  = NewRowY[212];
  assign \U52/DATA1_21  = NewRowY[213];
  assign \U52/DATA1_22  = NewRowY[214];
  assign \U52/DATA1_23  = NewRowY[215];
  assign \U52/DATA1_24  = NewRowY[216];
  assign \U52/DATA1_25  = NewRowY[217];
  assign \U52/DATA1_26  = NewRowY[218];
  assign \U52/DATA1_27  = NewRowY[219];
  assign \U52/DATA1_28  = NewRowY[220];
  assign \U52/DATA1_29  = NewRowY[221];
  assign \U52/DATA1_30  = NewRowY[222];
  assign \U52/DATA1_31  = NewRowY[223];
  assign \U52/DATA1_32  = NewRowY[224];
  assign \U52/DATA1_33  = NewRowY[225];
  assign \U52/DATA1_34  = NewRowY[226];
  assign \U52/DATA1_35  = NewRowY[227];
  assign \U52/DATA1_36  = NewRowY[228];
  assign \U52/DATA1_37  = NewRowY[229];
  assign \U52/DATA1_38  = NewRowY[230];
  assign \U52/DATA1_39  = NewRowY[231];
  assign \U52/DATA1_40  = NewRowY[232];
  assign \U52/DATA1_41  = NewRowY[233];
  assign \U52/DATA1_42  = NewRowY[234];
  assign \U52/DATA1_43  = NewRowY[235];
  assign \U52/DATA1_44  = NewRowY[236];
  assign \U52/DATA1_45  = NewRowY[237];
  assign \U52/DATA1_46  = NewRowY[238];
  assign \U52/DATA1_47  = NewRowY[239];
  assign \eq_207/A[15]  = NewRowY[255];
  assign \eq_207/A[14]  = NewRowY[254];
  assign \eq_207/A[13]  = NewRowY[253];
  assign \eq_207/A[12]  = NewRowY[252];
  assign \eq_207/A[11]  = NewRowY[251];
  assign \eq_207/A[10]  = NewRowY[250];
  assign \eq_207/A[9]  = NewRowY[249];
  assign \eq_207/A[8]  = NewRowY[248];
  assign \eq_207/A[7]  = NewRowY[247];
  assign \eq_207/A[6]  = NewRowY[246];
  assign \eq_207/A[5]  = NewRowY[245];
  assign \eq_207/A[4]  = NewRowY[244];
  assign \eq_207/A[3]  = NewRowY[243];
  assign \eq_207/A[2]  = NewRowY[242];
  assign \eq_207/A[1]  = NewRowY[241];
  assign \eq_207/A[0]  = NewRowY[240];
  assign \eq_207/B[15]  = X[15];
  assign \eq_207/B[14]  = X[14];
  assign \eq_207/B[13]  = X[13];
  assign \eq_207/B[12]  = X[12];
  assign \eq_207/B[11]  = X[11];
  assign \eq_207/B[10]  = X[10];
  assign \eq_207/B[9]  = X[9];
  assign \eq_207/B[8]  = X[8];
  assign \eq_207/B[7]  = X[7];
  assign \eq_207/B[6]  = X[6];
  assign \eq_207/B[5]  = X[5];
  assign \eq_207/B[4]  = X[4];
  assign \eq_207/B[3]  = X[3];
  assign \eq_207/B[2]  = X[2];
  assign \eq_207/B[1]  = X[1];
  assign \eq_207/B[0]  = X[0];
  assign \eq_112/A[15]  = NewRowX[255];
  assign \eq_112/A[14]  = NewRowX[254];
  assign \eq_112/A[13]  = NewRowX[253];
  assign \eq_112/A[12]  = NewRowX[252];
  assign \eq_112/A[11]  = NewRowX[251];
  assign \eq_112/A[10]  = NewRowX[250];
  assign \eq_112/A[9]  = NewRowX[249];
  assign \eq_112/A[8]  = NewRowX[248];
  assign \eq_112/A[7]  = NewRowX[247];
  assign \eq_112/A[6]  = NewRowX[246];
  assign \eq_112/A[5]  = NewRowX[245];
  assign \eq_112/A[4]  = NewRowX[244];
  assign \eq_112/A[3]  = NewRowX[243];
  assign \eq_112/A[2]  = NewRowX[242];
  assign \eq_112/A[1]  = NewRowX[241];
  assign \eq_112/A[0]  = NewRowX[240];
  assign \eq_112/B[15]  = Y[15];
  assign \eq_112/B[14]  = Y[14];
  assign \eq_112/B[13]  = Y[13];
  assign \eq_112/B[12]  = Y[12];
  assign \eq_112/B[11]  = Y[11];
  assign \eq_112/B[10]  = Y[10];
  assign \eq_112/B[9]  = Y[9];
  assign \eq_112/B[8]  = Y[8];
  assign \eq_112/B[7]  = Y[7];
  assign \eq_112/B[6]  = Y[6];
  assign \eq_112/B[5]  = Y[5];
  assign \eq_112/B[4]  = Y[4];
  assign \eq_112/B[3]  = Y[3];
  assign \eq_112/B[2]  = Y[2];
  assign \eq_112/B[1]  = Y[1];
  assign \eq_112/B[0]  = Y[0];
  assign \r528/A[15]  = NewRowY[63];
  assign \r528/A[14]  = NewRowY[62];
  assign \r528/A[13]  = NewRowY[61];
  assign \r528/A[12]  = NewRowY[60];
  assign \r528/A[11]  = NewRowY[59];
  assign \r528/A[10]  = NewRowY[58];
  assign \r528/A[9]  = NewRowY[57];
  assign \r528/A[8]  = NewRowY[56];
  assign \r528/A[7]  = NewRowY[55];
  assign \r528/A[6]  = NewRowY[54];
  assign \r528/A[5]  = NewRowY[53];
  assign \r528/A[4]  = NewRowY[52];
  assign \r528/A[3]  = NewRowY[51];
  assign \r528/A[2]  = NewRowY[50];
  assign \r528/A[1]  = NewRowY[49];
  assign \r528/A[0]  = NewRowY[48];
  assign \r527/A[15]  = NewRowY[127];
  assign \r527/A[14]  = NewRowY[126];
  assign \r527/A[13]  = NewRowY[125];
  assign \r527/A[12]  = NewRowY[124];
  assign \r527/A[11]  = NewRowY[123];
  assign \r527/A[10]  = NewRowY[122];
  assign \r527/A[9]  = NewRowY[121];
  assign \r527/A[8]  = NewRowY[120];
  assign \r527/A[7]  = NewRowY[119];
  assign \r527/A[6]  = NewRowY[118];
  assign \r527/A[5]  = NewRowY[117];
  assign \r527/A[4]  = NewRowY[116];
  assign \r527/A[3]  = NewRowY[115];
  assign \r527/A[2]  = NewRowY[114];
  assign \r527/A[1]  = NewRowY[113];
  assign \r527/A[0]  = NewRowY[112];
  assign \r526/A[15]  = NewRowY[191];
  assign \r526/A[14]  = NewRowY[190];
  assign \r526/A[13]  = NewRowY[189];
  assign \r526/A[12]  = NewRowY[188];
  assign \r526/A[11]  = NewRowY[187];
  assign \r526/A[10]  = NewRowY[186];
  assign \r526/A[9]  = NewRowY[185];
  assign \r526/A[8]  = NewRowY[184];
  assign \r526/A[7]  = NewRowY[183];
  assign \r526/A[6]  = NewRowY[182];
  assign \r526/A[5]  = NewRowY[181];
  assign \r526/A[4]  = NewRowY[180];
  assign \r526/A[3]  = NewRowY[179];
  assign \r526/A[2]  = NewRowY[178];
  assign \r526/A[1]  = NewRowY[177];
  assign \r526/A[0]  = NewRowY[176];
  assign \r524/A[15]  = NewRowX[63];
  assign \r524/A[14]  = NewRowX[62];
  assign \r524/A[13]  = NewRowX[61];
  assign \r524/A[12]  = NewRowX[60];
  assign \r524/A[11]  = NewRowX[59];
  assign \r524/A[10]  = NewRowX[58];
  assign \r524/A[9]  = NewRowX[57];
  assign \r524/A[8]  = NewRowX[56];
  assign \r524/A[7]  = NewRowX[55];
  assign \r524/A[6]  = NewRowX[54];
  assign \r524/A[5]  = NewRowX[53];
  assign \r524/A[4]  = NewRowX[52];
  assign \r524/A[3]  = NewRowX[51];
  assign \r524/A[2]  = NewRowX[50];
  assign \r524/A[1]  = NewRowX[49];
  assign \r524/A[0]  = NewRowX[48];
  assign \r523/A[15]  = NewRowX[127];
  assign \r523/A[14]  = NewRowX[126];
  assign \r523/A[13]  = NewRowX[125];
  assign \r523/A[12]  = NewRowX[124];
  assign \r523/A[11]  = NewRowX[123];
  assign \r523/A[10]  = NewRowX[122];
  assign \r523/A[9]  = NewRowX[121];
  assign \r523/A[8]  = NewRowX[120];
  assign \r523/A[7]  = NewRowX[119];
  assign \r523/A[6]  = NewRowX[118];
  assign \r523/A[5]  = NewRowX[117];
  assign \r523/A[4]  = NewRowX[116];
  assign \r523/A[3]  = NewRowX[115];
  assign \r523/A[2]  = NewRowX[114];
  assign \r523/A[1]  = NewRowX[113];
  assign \r523/A[0]  = NewRowX[112];
  assign \r522/A[15]  = NewRowX[191];
  assign \r522/A[14]  = NewRowX[190];
  assign \r522/A[13]  = NewRowX[189];
  assign \r522/A[12]  = NewRowX[188];
  assign \r522/A[11]  = NewRowX[187];
  assign \r522/A[10]  = NewRowX[186];
  assign \r522/A[9]  = NewRowX[185];
  assign \r522/A[8]  = NewRowX[184];
  assign \r522/A[7]  = NewRowX[183];
  assign \r522/A[6]  = NewRowX[182];
  assign \r522/A[5]  = NewRowX[181];
  assign \r522/A[4]  = NewRowX[180];
  assign \r522/A[3]  = NewRowX[179];
  assign \r522/A[2]  = NewRowX[178];
  assign \r522/A[1]  = NewRowX[177];
  assign \r522/A[0]  = NewRowX[176];

  DFF_X1 \FoundY_reg[0]  ( .D(n1078), .CK(clock), .Q(FoundY[0]), .QN(n29) );
  DFF_X1 \PosRowY_reg[1]  ( .D(n1075), .CK(clock), .Q(PosRowY[1]) );
  DFF_X1 \PosRowY_reg[0]  ( .D(n1076), .CK(clock), .Q(PosRowY[0]) );
  DFF_X1 \PosRowY_reg[2]  ( .D(n3928), .CK(clock), .Q(PosRowY[2]) );
  DFF_X1 \PosRowY_reg[3]  ( .D(n3929), .CK(clock), .Q(PosRowY[3]) );
  DFF_X1 \PosRowY_reg[4]  ( .D(n3930), .CK(clock), .Q(PosRowY[4]) );
  DFF_X1 \PosRowY_reg[5]  ( .D(n3931), .CK(clock), .Q(PosRowY[5]) );
  DFF_X1 \PosRowY_reg[6]  ( .D(n3932), .CK(clock), .Q(PosRowY[6]) );
  DFF_X1 \PosRowY_reg[7]  ( .D(n3933), .CK(clock), .Q(PosRowY[7]) );
  DFF_X1 \PosRowY_reg[8]  ( .D(n3934), .CK(clock), .Q(PosRowY[8]) );
  DFF_X1 \PosRowY_reg[9]  ( .D(n3935), .CK(clock), .Q(PosRowY[9]) );
  DFF_X1 \PosRowY_reg[10]  ( .D(n3936), .CK(clock), .Q(PosRowY[10]) );
  DFF_X1 \PosRowY_reg[11]  ( .D(n3937), .CK(clock), .Q(PosRowY[11]) );
  DFF_X1 \PosRowY_reg[12]  ( .D(n3938), .CK(clock), .Q(PosRowY[12]) );
  DFF_X1 \FoundX_reg[0]  ( .D(n1074), .CK(clock), .Q(FoundX[0]), .QN(n36) );
  DFF_X1 \PosRowX_reg[1]  ( .D(n1023), .CK(clock), .Q(PosRowX[1]) );
  DFF_X1 \PosRowX_reg[0]  ( .D(n1024), .CK(clock), .Q(PosRowX[0]) );
  DFF_X1 \PosRowX_reg[2]  ( .D(n3942), .CK(clock), .Q(PosRowX[2]) );
  DFF_X1 \PosRowX_reg[3]  ( .D(n3943), .CK(clock), .Q(PosRowX[3]) );
  DFF_X1 \PosRowX_reg[4]  ( .D(n3944), .CK(clock), .Q(PosRowX[4]) );
  DFF_X1 \PosRowX_reg[5]  ( .D(n3945), .CK(clock), .Q(PosRowX[5]) );
  DFF_X1 \PosRowX_reg[6]  ( .D(n3946), .CK(clock), .Q(PosRowX[6]) );
  DFF_X1 \PosRowX_reg[7]  ( .D(n3947), .CK(clock), .Q(PosRowX[7]) );
  DFF_X1 \PosRowX_reg[8]  ( .D(n3948), .CK(clock), .Q(PosRowX[8]) );
  DFF_X1 \PosRowX_reg[9]  ( .D(n3949), .CK(clock), .Q(PosRowX[9]) );
  DFF_X1 \PosRowX_reg[10]  ( .D(n3950), .CK(clock), .Q(PosRowX[10]) );
  DFF_X1 \PosRowX_reg[11]  ( .D(n3951), .CK(clock), .Q(PosRowX[11]) );
  DFF_X1 \PosRowX_reg[12]  ( .D(n3952), .CK(clock), .Q(PosRowX[12]) );
  DFF_X1 \Element_reg[47]  ( .D(n1025), .CK(clock), .Q(Element[47]) );
  DFF_X1 \Element_reg[46]  ( .D(n1026), .CK(clock), .Q(Element[46]) );
  DFF_X1 \Element_reg[45]  ( .D(n1027), .CK(clock), .Q(Element[45]) );
  DFF_X1 \Element_reg[44]  ( .D(n1028), .CK(clock), .Q(Element[44]) );
  DFF_X1 \Element_reg[43]  ( .D(n1029), .CK(clock), .Q(Element[43]) );
  DFF_X1 \Element_reg[42]  ( .D(n1030), .CK(clock), .Q(Element[42]) );
  DFF_X1 \Element_reg[41]  ( .D(n1031), .CK(clock), .Q(Element[41]) );
  DFF_X1 \Element_reg[40]  ( .D(n1032), .CK(clock), .Q(Element[40]) );
  DFF_X1 \Element_reg[39]  ( .D(n1033), .CK(clock), .Q(Element[39]) );
  DFF_X1 \Element_reg[38]  ( .D(n1034), .CK(clock), .Q(Element[38]) );
  DFF_X1 \Element_reg[37]  ( .D(n1035), .CK(clock), .Q(Element[37]) );
  DFF_X1 \Element_reg[36]  ( .D(n1036), .CK(clock), .Q(Element[36]) );
  DFF_X1 \Element_reg[35]  ( .D(n1037), .CK(clock), .Q(Element[35]) );
  DFF_X1 \Element_reg[34]  ( .D(n1038), .CK(clock), .Q(Element[34]) );
  DFF_X1 \Element_reg[33]  ( .D(n1039), .CK(clock), .Q(Element[33]) );
  DFF_X1 \Element_reg[32]  ( .D(n1040), .CK(clock), .Q(Element[32]) );
  DFF_X1 \Element_reg[31]  ( .D(n1041), .CK(clock), .Q(Element[31]) );
  DFF_X1 \Element_reg[30]  ( .D(n1042), .CK(clock), .Q(Element[30]) );
  DFF_X1 \Element_reg[29]  ( .D(n1043), .CK(clock), .Q(Element[29]) );
  DFF_X1 \Element_reg[28]  ( .D(n1044), .CK(clock), .Q(Element[28]) );
  DFF_X1 \Element_reg[27]  ( .D(n1045), .CK(clock), .Q(Element[27]) );
  DFF_X1 \Element_reg[26]  ( .D(n1046), .CK(clock), .Q(Element[26]) );
  DFF_X1 \Element_reg[25]  ( .D(n1047), .CK(clock), .Q(Element[25]) );
  DFF_X1 \Element_reg[24]  ( .D(n1048), .CK(clock), .Q(Element[24]) );
  DFF_X1 \Element_reg[23]  ( .D(n1049), .CK(clock), .Q(Element[23]) );
  DFF_X1 \Element_reg[22]  ( .D(n1050), .CK(clock), .Q(Element[22]) );
  DFF_X1 \Element_reg[21]  ( .D(n1051), .CK(clock), .Q(Element[21]) );
  DFF_X1 \Element_reg[20]  ( .D(n1052), .CK(clock), .Q(Element[20]) );
  DFF_X1 \Element_reg[19]  ( .D(n1053), .CK(clock), .Q(Element[19]) );
  DFF_X1 \Element_reg[18]  ( .D(n1054), .CK(clock), .Q(Element[18]) );
  DFF_X1 \Element_reg[17]  ( .D(n1055), .CK(clock), .Q(Element[17]) );
  DFF_X1 \Element_reg[16]  ( .D(n1056), .CK(clock), .Q(Element[16]) );
  DFF_X1 \Element_reg[15]  ( .D(n1057), .CK(clock), .Q(Element[15]) );
  DFF_X1 \Element_reg[14]  ( .D(n1058), .CK(clock), .Q(Element[14]) );
  DFF_X1 \Element_reg[13]  ( .D(n1059), .CK(clock), .Q(Element[13]) );
  DFF_X1 \Element_reg[12]  ( .D(n1060), .CK(clock), .Q(Element[12]) );
  DFF_X1 \Element_reg[11]  ( .D(n1061), .CK(clock), .Q(Element[11]) );
  DFF_X1 \Element_reg[10]  ( .D(n1062), .CK(clock), .Q(Element[10]) );
  DFF_X1 \Element_reg[9]  ( .D(n1063), .CK(clock), .Q(Element[9]) );
  DFF_X1 \Element_reg[8]  ( .D(n1064), .CK(clock), .Q(Element[8]) );
  DFF_X1 \Element_reg[7]  ( .D(n1065), .CK(clock), .Q(Element[7]) );
  DFF_X1 \Element_reg[6]  ( .D(n1066), .CK(clock), .Q(Element[6]) );
  DFF_X1 \Element_reg[5]  ( .D(n1067), .CK(clock), .Q(Element[5]) );
  DFF_X1 \Element_reg[4]  ( .D(n1068), .CK(clock), .Q(Element[4]) );
  DFF_X1 \Element_reg[3]  ( .D(n1069), .CK(clock), .Q(Element[3]) );
  DFF_X1 \Element_reg[2]  ( .D(n1070), .CK(clock), .Q(Element[2]) );
  DFF_X1 \Element_reg[1]  ( .D(n1071), .CK(clock), .Q(Element[1]) );
  DFF_X1 \Element_reg[0]  ( .D(n1072), .CK(clock), .Q(Element[0]) );
  NAND2_X2 U4 ( .A1(PosRowX[1]), .A2(n3953), .ZN(n194) );
  OAI221_X2 U7 ( .B1(n197), .B2(n3954), .C1(n198), .C2(n3966), .A(n3926), .ZN(
        n196) );
  OAI221_X2 U23 ( .B1(n4063), .B2(n226), .C1(n221), .C2(n3893), .A(n228), .ZN(
        n223) );
  AOI221_X2 U25 ( .B1(n3914), .B2(\U168/DATA1_47 ), .C1(n3940), .C2(n234), .A(
        n235), .ZN(n232) );
  OAI221_X2 U27 ( .B1(n3967), .B2(n3899), .C1(n4015), .C2(n3897), .A(n239), 
        .ZN(n234) );
  OAI221_X2 U35 ( .B1(n3916), .B2(n4064), .C1(n3893), .C2(n251), .A(n253), 
        .ZN(n252) );
  AOI221_X2 U37 ( .B1(\U168/DATA1_46 ), .B2(n3914), .C1(n3910), .C2(n256), .A(
        n257), .ZN(n255) );
  OAI221_X2 U39 ( .B1(n3899), .B2(n3968), .C1(n3897), .C2(n4016), .A(n258), 
        .ZN(n256) );
  OAI221_X2 U47 ( .B1(n226), .B2(n4065), .C1(n3893), .C2(n263), .A(n265), .ZN(
        n264) );
  AOI221_X2 U49 ( .B1(\U168/DATA1_45 ), .B2(n3913), .C1(n3910), .C2(n268), .A(
        n269), .ZN(n267) );
  OAI221_X2 U51 ( .B1(n3899), .B2(n3969), .C1(n3897), .C2(n4017), .A(n270), 
        .ZN(n268) );
  OAI221_X2 U59 ( .B1(n3916), .B2(n4066), .C1(n3893), .C2(n275), .A(n277), 
        .ZN(n276) );
  AOI221_X2 U61 ( .B1(\U168/DATA1_44 ), .B2(n3913), .C1(n3910), .C2(n280), .A(
        n281), .ZN(n279) );
  OAI221_X2 U63 ( .B1(n3899), .B2(n3970), .C1(n3897), .C2(n4018), .A(n282), 
        .ZN(n280) );
  OAI221_X2 U71 ( .B1(n226), .B2(n4067), .C1(n3893), .C2(n287), .A(n289), .ZN(
        n288) );
  AOI221_X2 U73 ( .B1(\U168/DATA1_43 ), .B2(n3914), .C1(n3940), .C2(n292), .A(
        n293), .ZN(n291) );
  OAI221_X2 U75 ( .B1(n3899), .B2(n3971), .C1(n3897), .C2(n4019), .A(n294), 
        .ZN(n292) );
  OAI221_X2 U83 ( .B1(n3916), .B2(n4068), .C1(n3893), .C2(n299), .A(n301), 
        .ZN(n300) );
  AOI221_X2 U85 ( .B1(\U168/DATA1_42 ), .B2(n3914), .C1(n3910), .C2(n304), .A(
        n305), .ZN(n303) );
  OAI221_X2 U87 ( .B1(n3899), .B2(n3972), .C1(n3897), .C2(n4020), .A(n306), 
        .ZN(n304) );
  OAI221_X2 U95 ( .B1(n226), .B2(n4069), .C1(n3893), .C2(n311), .A(n313), .ZN(
        n312) );
  AOI221_X2 U97 ( .B1(\U168/DATA1_41 ), .B2(n3913), .C1(n3910), .C2(n316), .A(
        n317), .ZN(n315) );
  OAI221_X2 U99 ( .B1(n3899), .B2(n3973), .C1(n3897), .C2(n4021), .A(n318), 
        .ZN(n316) );
  OAI221_X2 U107 ( .B1(n226), .B2(n4070), .C1(n3893), .C2(n323), .A(n325), 
        .ZN(n324) );
  AOI221_X2 U109 ( .B1(\U168/DATA1_40 ), .B2(n3914), .C1(n3910), .C2(n328), 
        .A(n329), .ZN(n327) );
  OAI221_X2 U111 ( .B1(n3899), .B2(n3974), .C1(n3897), .C2(n4022), .A(n330), 
        .ZN(n328) );
  OAI221_X2 U119 ( .B1(n226), .B2(n4071), .C1(n3893), .C2(n335), .A(n337), 
        .ZN(n336) );
  AOI221_X2 U121 ( .B1(\U168/DATA1_39 ), .B2(n3913), .C1(n3940), .C2(n340), 
        .A(n341), .ZN(n339) );
  OAI221_X2 U123 ( .B1(n3899), .B2(n3975), .C1(n3897), .C2(n4023), .A(n342), 
        .ZN(n340) );
  OAI221_X2 U131 ( .B1(n226), .B2(n4072), .C1(n3893), .C2(n347), .A(n349), 
        .ZN(n348) );
  AOI221_X2 U133 ( .B1(\U168/DATA1_38 ), .B2(n3914), .C1(n3910), .C2(n352), 
        .A(n353), .ZN(n351) );
  OAI221_X2 U135 ( .B1(n3899), .B2(n3976), .C1(n3897), .C2(n4024), .A(n354), 
        .ZN(n352) );
  OAI221_X2 U143 ( .B1(n226), .B2(n4073), .C1(n3893), .C2(n359), .A(n361), 
        .ZN(n360) );
  AOI221_X2 U145 ( .B1(\U168/DATA1_37 ), .B2(n3914), .C1(n3910), .C2(n364), 
        .A(n365), .ZN(n363) );
  OAI221_X2 U147 ( .B1(n3899), .B2(n3977), .C1(n3897), .C2(n4025), .A(n366), 
        .ZN(n364) );
  OAI221_X2 U155 ( .B1(n226), .B2(n4074), .C1(n3893), .C2(n371), .A(n373), 
        .ZN(n372) );
  AOI221_X2 U157 ( .B1(\U168/DATA1_36 ), .B2(n3914), .C1(n3940), .C2(n376), 
        .A(n377), .ZN(n375) );
  OAI221_X2 U159 ( .B1(n3899), .B2(n3978), .C1(n3897), .C2(n4026), .A(n378), 
        .ZN(n376) );
  OAI221_X2 U167 ( .B1(n226), .B2(n4075), .C1(n3893), .C2(n383), .A(n385), 
        .ZN(n384) );
  AOI221_X2 U169 ( .B1(\U168/DATA1_35 ), .B2(n3914), .C1(n3910), .C2(n388), 
        .A(n389), .ZN(n387) );
  OAI221_X2 U171 ( .B1(n3899), .B2(n3979), .C1(n3897), .C2(n4027), .A(n390), 
        .ZN(n388) );
  OAI221_X2 U179 ( .B1(n3916), .B2(n4076), .C1(n3893), .C2(n395), .A(n397), 
        .ZN(n396) );
  AOI221_X2 U181 ( .B1(\U168/DATA1_34 ), .B2(n3914), .C1(n3940), .C2(n400), 
        .A(n401), .ZN(n399) );
  OAI221_X2 U183 ( .B1(n3899), .B2(n3980), .C1(n3897), .C2(n4028), .A(n402), 
        .ZN(n400) );
  OAI221_X2 U191 ( .B1(n3916), .B2(n4077), .C1(n3893), .C2(n407), .A(n409), 
        .ZN(n408) );
  AOI221_X2 U193 ( .B1(\U168/DATA1_33 ), .B2(n3914), .C1(n3910), .C2(n412), 
        .A(n413), .ZN(n411) );
  OAI221_X2 U195 ( .B1(n3899), .B2(n3981), .C1(n3897), .C2(n4029), .A(n414), 
        .ZN(n412) );
  OAI221_X2 U203 ( .B1(n3916), .B2(n4078), .C1(n3893), .C2(n419), .A(n421), 
        .ZN(n420) );
  AOI221_X2 U205 ( .B1(\U168/DATA1_32 ), .B2(n3914), .C1(n3940), .C2(n424), 
        .A(n425), .ZN(n423) );
  OAI221_X2 U207 ( .B1(n3899), .B2(n3982), .C1(n3897), .C2(n4030), .A(n426), 
        .ZN(n424) );
  OAI221_X2 U215 ( .B1(n3916), .B2(n4079), .C1(n3893), .C2(n431), .A(n433), 
        .ZN(n432) );
  AOI221_X2 U217 ( .B1(\U168/DATA1_31 ), .B2(n3914), .C1(n3910), .C2(n436), 
        .A(n437), .ZN(n435) );
  OAI221_X2 U219 ( .B1(n3899), .B2(n3983), .C1(n3897), .C2(n4031), .A(n438), 
        .ZN(n436) );
  OAI221_X2 U227 ( .B1(n3916), .B2(n4080), .C1(n3893), .C2(n443), .A(n445), 
        .ZN(n444) );
  AOI221_X2 U229 ( .B1(\U168/DATA1_30 ), .B2(n3914), .C1(n3940), .C2(n448), 
        .A(n449), .ZN(n447) );
  OAI221_X2 U231 ( .B1(n3899), .B2(n3984), .C1(n3897), .C2(n4032), .A(n450), 
        .ZN(n448) );
  OAI221_X2 U239 ( .B1(n3916), .B2(n4081), .C1(n3893), .C2(n455), .A(n457), 
        .ZN(n456) );
  AOI221_X2 U241 ( .B1(\U168/DATA1_29 ), .B2(n3914), .C1(n3910), .C2(n460), 
        .A(n461), .ZN(n459) );
  OAI221_X2 U243 ( .B1(n3899), .B2(n3985), .C1(n3897), .C2(n4033), .A(n462), 
        .ZN(n460) );
  OAI221_X2 U251 ( .B1(n3916), .B2(n4082), .C1(n3893), .C2(n467), .A(n469), 
        .ZN(n468) );
  AOI221_X2 U253 ( .B1(\U168/DATA1_28 ), .B2(n3914), .C1(n3910), .C2(n472), 
        .A(n473), .ZN(n471) );
  OAI221_X2 U255 ( .B1(n3899), .B2(n3986), .C1(n3897), .C2(n4034), .A(n474), 
        .ZN(n472) );
  OAI221_X2 U263 ( .B1(n3916), .B2(n4083), .C1(n3893), .C2(n479), .A(n481), 
        .ZN(n480) );
  AOI221_X2 U265 ( .B1(\U168/DATA1_27 ), .B2(n3914), .C1(n3940), .C2(n484), 
        .A(n485), .ZN(n483) );
  OAI221_X2 U267 ( .B1(n3899), .B2(n3987), .C1(n3897), .C2(n4035), .A(n486), 
        .ZN(n484) );
  OAI221_X2 U275 ( .B1(n3916), .B2(n4084), .C1(n3893), .C2(n491), .A(n493), 
        .ZN(n492) );
  AOI221_X2 U277 ( .B1(\U168/DATA1_26 ), .B2(n3914), .C1(n3910), .C2(n496), 
        .A(n497), .ZN(n495) );
  OAI221_X2 U279 ( .B1(n3899), .B2(n3988), .C1(n3897), .C2(n4036), .A(n498), 
        .ZN(n496) );
  OAI221_X2 U287 ( .B1(n3916), .B2(n4085), .C1(n3893), .C2(n503), .A(n505), 
        .ZN(n504) );
  AOI221_X2 U289 ( .B1(\U168/DATA1_25 ), .B2(n3913), .C1(n3910), .C2(n508), 
        .A(n509), .ZN(n507) );
  OAI221_X2 U291 ( .B1(n3899), .B2(n3989), .C1(n3897), .C2(n4037), .A(n510), 
        .ZN(n508) );
  OAI221_X2 U299 ( .B1(n3916), .B2(n4086), .C1(n3893), .C2(n515), .A(n517), 
        .ZN(n516) );
  AOI221_X2 U301 ( .B1(\U168/DATA1_24 ), .B2(n3913), .C1(n3910), .C2(n520), 
        .A(n521), .ZN(n519) );
  OAI221_X2 U303 ( .B1(n3899), .B2(n3990), .C1(n3897), .C2(n4038), .A(n522), 
        .ZN(n520) );
  OAI221_X2 U311 ( .B1(n3916), .B2(n4087), .C1(n3893), .C2(n527), .A(n529), 
        .ZN(n528) );
  AOI221_X2 U313 ( .B1(\U168/DATA1_23 ), .B2(n3913), .C1(n3910), .C2(n532), 
        .A(n533), .ZN(n531) );
  OAI221_X2 U315 ( .B1(n3899), .B2(n3991), .C1(n3897), .C2(n4039), .A(n534), 
        .ZN(n532) );
  OAI221_X2 U323 ( .B1(n3916), .B2(n4088), .C1(n3893), .C2(n539), .A(n541), 
        .ZN(n540) );
  AOI221_X2 U325 ( .B1(\U168/DATA1_22 ), .B2(n3913), .C1(n3910), .C2(n544), 
        .A(n545), .ZN(n543) );
  OAI221_X2 U327 ( .B1(n3899), .B2(n3992), .C1(n3897), .C2(n4040), .A(n546), 
        .ZN(n544) );
  OAI221_X2 U335 ( .B1(n226), .B2(n4089), .C1(n3893), .C2(n551), .A(n553), 
        .ZN(n552) );
  AOI221_X2 U337 ( .B1(\U168/DATA1_21 ), .B2(n3913), .C1(n3910), .C2(n556), 
        .A(n557), .ZN(n555) );
  OAI221_X2 U339 ( .B1(n3899), .B2(n3993), .C1(n3897), .C2(n4041), .A(n558), 
        .ZN(n556) );
  OAI221_X2 U347 ( .B1(n226), .B2(n4090), .C1(n3893), .C2(n563), .A(n565), 
        .ZN(n564) );
  AOI221_X2 U349 ( .B1(\U168/DATA1_20 ), .B2(n3913), .C1(n3910), .C2(n568), 
        .A(n569), .ZN(n567) );
  OAI221_X2 U351 ( .B1(n3899), .B2(n3994), .C1(n3897), .C2(n4042), .A(n570), 
        .ZN(n568) );
  OAI221_X2 U359 ( .B1(n226), .B2(n4091), .C1(n3893), .C2(n575), .A(n577), 
        .ZN(n576) );
  AOI221_X2 U361 ( .B1(\U168/DATA1_19 ), .B2(n3913), .C1(n3910), .C2(n580), 
        .A(n581), .ZN(n579) );
  OAI221_X2 U363 ( .B1(n3899), .B2(n3995), .C1(n3897), .C2(n4043), .A(n582), 
        .ZN(n580) );
  OAI221_X2 U371 ( .B1(n226), .B2(n4092), .C1(n3893), .C2(n587), .A(n589), 
        .ZN(n588) );
  AOI221_X2 U373 ( .B1(\U168/DATA1_18 ), .B2(n3913), .C1(n3910), .C2(n592), 
        .A(n593), .ZN(n591) );
  OAI221_X2 U375 ( .B1(n3899), .B2(n3996), .C1(n3897), .C2(n4044), .A(n594), 
        .ZN(n592) );
  OAI221_X2 U383 ( .B1(n226), .B2(n4093), .C1(n3893), .C2(n599), .A(n601), 
        .ZN(n600) );
  AOI221_X2 U385 ( .B1(\U168/DATA1_17 ), .B2(n3913), .C1(n3910), .C2(n604), 
        .A(n605), .ZN(n603) );
  OAI221_X2 U387 ( .B1(n3899), .B2(n3997), .C1(n3897), .C2(n4045), .A(n606), 
        .ZN(n604) );
  OAI221_X2 U395 ( .B1(n226), .B2(n4094), .C1(n3893), .C2(n611), .A(n613), 
        .ZN(n612) );
  AOI221_X2 U397 ( .B1(\U168/DATA1_16 ), .B2(n3913), .C1(n3910), .C2(n616), 
        .A(n617), .ZN(n615) );
  OAI221_X2 U399 ( .B1(n3899), .B2(n3998), .C1(n3897), .C2(n4046), .A(n618), 
        .ZN(n616) );
  OAI221_X2 U407 ( .B1(n226), .B2(n4095), .C1(n3893), .C2(n623), .A(n625), 
        .ZN(n624) );
  AOI221_X2 U409 ( .B1(\U168/DATA1_15 ), .B2(n3913), .C1(n3910), .C2(n628), 
        .A(n629), .ZN(n627) );
  OAI221_X2 U411 ( .B1(n3899), .B2(n3999), .C1(n3897), .C2(n4047), .A(n630), 
        .ZN(n628) );
  OAI221_X2 U419 ( .B1(n3916), .B2(n4096), .C1(n3893), .C2(n635), .A(n637), 
        .ZN(n636) );
  AOI221_X2 U421 ( .B1(\U168/DATA1_14 ), .B2(n3913), .C1(n3910), .C2(n640), 
        .A(n641), .ZN(n639) );
  OAI221_X2 U423 ( .B1(n3899), .B2(n4000), .C1(n3897), .C2(n4048), .A(n642), 
        .ZN(n640) );
  OAI221_X2 U431 ( .B1(n3916), .B2(n4097), .C1(n3893), .C2(n647), .A(n649), 
        .ZN(n648) );
  AOI221_X2 U433 ( .B1(\U168/DATA1_13 ), .B2(n3913), .C1(n3910), .C2(n652), 
        .A(n653), .ZN(n651) );
  OAI221_X2 U435 ( .B1(n3899), .B2(n4001), .C1(n3897), .C2(n4049), .A(n654), 
        .ZN(n652) );
  OAI221_X2 U443 ( .B1(n226), .B2(n4098), .C1(n3893), .C2(n659), .A(n661), 
        .ZN(n660) );
  AOI221_X2 U445 ( .B1(\U168/DATA1_12 ), .B2(n3913), .C1(n3940), .C2(n664), 
        .A(n665), .ZN(n663) );
  OAI221_X2 U447 ( .B1(n3899), .B2(n4002), .C1(n3897), .C2(n4050), .A(n666), 
        .ZN(n664) );
  OAI221_X2 U455 ( .B1(n3916), .B2(n4099), .C1(n3893), .C2(n671), .A(n673), 
        .ZN(n672) );
  AOI221_X2 U457 ( .B1(\U168/DATA1_11 ), .B2(n3914), .C1(n3940), .C2(n676), 
        .A(n677), .ZN(n675) );
  OAI221_X2 U459 ( .B1(n3899), .B2(n4003), .C1(n3897), .C2(n4051), .A(n678), 
        .ZN(n676) );
  OAI221_X2 U467 ( .B1(n3916), .B2(n4100), .C1(n3893), .C2(n683), .A(n685), 
        .ZN(n684) );
  AOI221_X2 U469 ( .B1(\U168/DATA1_10 ), .B2(n3914), .C1(n3940), .C2(n688), 
        .A(n689), .ZN(n687) );
  OAI221_X2 U471 ( .B1(n3899), .B2(n4004), .C1(n3897), .C2(n4052), .A(n690), 
        .ZN(n688) );
  OAI221_X2 U479 ( .B1(n3916), .B2(n4101), .C1(n3893), .C2(n695), .A(n697), 
        .ZN(n696) );
  AOI221_X2 U481 ( .B1(\U168/DATA1_9 ), .B2(n3913), .C1(n3940), .C2(n700), .A(
        n701), .ZN(n699) );
  OAI221_X2 U483 ( .B1(n3899), .B2(n4005), .C1(n3897), .C2(n4053), .A(n702), 
        .ZN(n700) );
  OAI221_X2 U491 ( .B1(n3916), .B2(n4102), .C1(n3893), .C2(n707), .A(n709), 
        .ZN(n708) );
  AOI221_X2 U493 ( .B1(\U168/DATA1_8 ), .B2(n3914), .C1(n3940), .C2(n712), .A(
        n713), .ZN(n711) );
  OAI221_X2 U495 ( .B1(n3899), .B2(n4006), .C1(n3897), .C2(n4054), .A(n714), 
        .ZN(n712) );
  OAI221_X2 U503 ( .B1(n226), .B2(n4103), .C1(n3893), .C2(n719), .A(n721), 
        .ZN(n720) );
  AOI221_X2 U505 ( .B1(\U168/DATA1_7 ), .B2(n3914), .C1(n3910), .C2(n724), .A(
        n725), .ZN(n723) );
  OAI221_X2 U507 ( .B1(n3899), .B2(n4007), .C1(n3897), .C2(n4055), .A(n726), 
        .ZN(n724) );
  OAI221_X2 U515 ( .B1(n3916), .B2(n4104), .C1(n3893), .C2(n731), .A(n733), 
        .ZN(n732) );
  AOI221_X2 U517 ( .B1(\U168/DATA1_6 ), .B2(n3913), .C1(n3940), .C2(n736), .A(
        n737), .ZN(n735) );
  OAI221_X2 U519 ( .B1(n3899), .B2(n4008), .C1(n3897), .C2(n4056), .A(n738), 
        .ZN(n736) );
  OAI221_X2 U527 ( .B1(n226), .B2(n4105), .C1(n3893), .C2(n743), .A(n745), 
        .ZN(n744) );
  AOI221_X2 U529 ( .B1(\U168/DATA1_5 ), .B2(n3913), .C1(n3910), .C2(n748), .A(
        n749), .ZN(n747) );
  OAI221_X2 U531 ( .B1(n3899), .B2(n4009), .C1(n3897), .C2(n4057), .A(n750), 
        .ZN(n748) );
  OAI221_X2 U539 ( .B1(n3916), .B2(n4106), .C1(n3893), .C2(n755), .A(n757), 
        .ZN(n756) );
  AOI221_X2 U541 ( .B1(\U168/DATA1_4 ), .B2(n3914), .C1(n3910), .C2(n760), .A(
        n761), .ZN(n759) );
  OAI221_X2 U543 ( .B1(n3899), .B2(n4010), .C1(n3897), .C2(n4058), .A(n762), 
        .ZN(n760) );
  OAI221_X2 U551 ( .B1(n226), .B2(n4107), .C1(n3893), .C2(n767), .A(n769), 
        .ZN(n768) );
  AOI221_X2 U553 ( .B1(\U168/DATA1_3 ), .B2(n3913), .C1(n3910), .C2(n772), .A(
        n773), .ZN(n771) );
  OAI221_X2 U555 ( .B1(n3899), .B2(n4011), .C1(n3897), .C2(n4059), .A(n774), 
        .ZN(n772) );
  OAI221_X2 U563 ( .B1(n3916), .B2(n4108), .C1(n3893), .C2(n779), .A(n781), 
        .ZN(n780) );
  AOI221_X2 U565 ( .B1(\U168/DATA1_2 ), .B2(n3913), .C1(n3910), .C2(n784), .A(
        n785), .ZN(n783) );
  OAI221_X2 U567 ( .B1(n3899), .B2(n4012), .C1(n3897), .C2(n4060), .A(n786), 
        .ZN(n784) );
  OAI221_X2 U575 ( .B1(n226), .B2(n4109), .C1(n3893), .C2(n791), .A(n793), 
        .ZN(n792) );
  AOI221_X2 U577 ( .B1(\U168/DATA1_1 ), .B2(n3914), .C1(n3910), .C2(n796), .A(
        n797), .ZN(n795) );
  OAI221_X2 U579 ( .B1(n3899), .B2(n4013), .C1(n3897), .C2(n4061), .A(n798), 
        .ZN(n796) );
  NAND2_X2 U587 ( .A1(n805), .A2(n3961), .ZN(n222) );
  OAI221_X2 U588 ( .B1(n3916), .B2(n4110), .C1(n3893), .C2(n803), .A(n806), 
        .ZN(n804) );
  AOI221_X2 U590 ( .B1(\U168/DATA1_0 ), .B2(n3913), .C1(n3940), .C2(n811), .A(
        n812), .ZN(n810) );
  OAI221_X2 U593 ( .B1(n3899), .B2(n4014), .C1(n3897), .C2(n4062), .A(n814), 
        .ZN(n811) );
  NOR2_X2 U597 ( .A1(n198), .A2(n3965), .ZN(n816) );
  NOR2_X2 U600 ( .A1(n822), .A2(n813), .ZN(n197) );
  NAND2_X2 U601 ( .A1(n807), .A2(n3963), .ZN(n226) );
  NOR3_X2 U602 ( .A1(n826), .A2(n827), .A3(n823), .ZN(n215) );
  NAND4_X2 U603 ( .A1(n828), .A2(n3896), .A3(n829), .A4(n830), .ZN(n824) );
  NAND2_X2 U605 ( .A1(n3955), .A2(WireX), .ZN(n829) );
  NOR2_X2 U608 ( .A1(n834), .A2(n3961), .ZN(n808) );
  OAI22_X2 U611 ( .A1(n36), .A2(n835), .B1(n3955), .B2(n818), .ZN(n1074) );
  NAND2_X2 U612 ( .A1(WireX), .A2(n838), .ZN(n818) );
  NAND3_X2 U613 ( .A1(n813), .A2(n3956), .A3(PosDX[1]), .ZN(n838) );
  NOR2_X2 U615 ( .A1(n3956), .A2(PosDX[1]), .ZN(n817) );
  NOR2_X2 U616 ( .A1(PosDX[1]), .A2(PosDX[0]), .ZN(n815) );
  NAND2_X2 U617 ( .A1(n832), .A2(n828), .ZN(n835) );
  NAND3_X2 U619 ( .A1(DiagonalDoneX), .A2(n35), .A3(FoundX[0]), .ZN(n819) );
  NAND2_X2 U620 ( .A1(n193), .A2(n198), .ZN(n820) );
  NAND4_X2 U621 ( .A1(n840), .A2(n841), .A3(n842), .A4(n843), .ZN(n198) );
  NOR4_X2 U622 ( .A1(n844), .A2(n845), .A3(n846), .A4(n847), .ZN(n843) );
  XOR2_X2 U623 ( .A(\r522/A[3] ), .B(\eq_112/B[3] ), .Z(n847) );
  XOR2_X2 U624 ( .A(\r522/A[2] ), .B(\eq_112/B[2] ), .Z(n846) );
  XOR2_X2 U625 ( .A(\r522/A[1] ), .B(\eq_112/B[1] ), .Z(n845) );
  XOR2_X2 U626 ( .A(\r522/A[0] ), .B(\eq_112/B[0] ), .Z(n844) );
  NOR4_X2 U627 ( .A1(n848), .A2(n849), .A3(n850), .A4(n851), .ZN(n842) );
  XOR2_X2 U628 ( .A(\r522/A[7] ), .B(\eq_112/B[7] ), .Z(n851) );
  XOR2_X2 U629 ( .A(\r522/A[6] ), .B(\eq_112/B[6] ), .Z(n850) );
  XOR2_X2 U630 ( .A(\r522/A[5] ), .B(\eq_112/B[5] ), .Z(n849) );
  XOR2_X2 U631 ( .A(\r522/A[4] ), .B(\eq_112/B[4] ), .Z(n848) );
  NOR4_X2 U632 ( .A1(n852), .A2(n853), .A3(n854), .A4(n855), .ZN(n841) );
  XOR2_X2 U633 ( .A(\r522/A[11] ), .B(\eq_112/B[11] ), .Z(n855) );
  XOR2_X2 U634 ( .A(\r522/A[10] ), .B(\eq_112/B[10] ), .Z(n854) );
  XOR2_X2 U635 ( .A(\r522/A[9] ), .B(\eq_112/B[9] ), .Z(n853) );
  XOR2_X2 U636 ( .A(\r522/A[8] ), .B(\eq_112/B[8] ), .Z(n852) );
  NOR4_X2 U637 ( .A1(n856), .A2(n857), .A3(n858), .A4(n859), .ZN(n840) );
  XOR2_X2 U638 ( .A(\r522/A[15] ), .B(\eq_112/B[15] ), .Z(n859) );
  XOR2_X2 U639 ( .A(\r522/A[14] ), .B(\eq_112/B[14] ), .Z(n858) );
  XOR2_X2 U640 ( .A(\r522/A[13] ), .B(\eq_112/B[13] ), .Z(n857) );
  XOR2_X2 U641 ( .A(\r522/A[12] ), .B(\eq_112/B[12] ), .Z(n856) );
  NOR2_X2 U642 ( .A1(n3966), .A2(n813), .ZN(n193) );
  AND4_X2 U643 ( .A1(n860), .A2(n861), .A3(n862), .A4(n863), .ZN(n813) );
  NOR4_X2 U644 ( .A1(n864), .A2(n865), .A3(n866), .A4(n867), .ZN(n863) );
  XOR2_X2 U645 ( .A(\r524/A[3] ), .B(\eq_112/B[3] ), .Z(n867) );
  XOR2_X2 U646 ( .A(\r524/A[2] ), .B(\eq_112/B[2] ), .Z(n866) );
  XOR2_X2 U647 ( .A(\r524/A[1] ), .B(\eq_112/B[1] ), .Z(n865) );
  XOR2_X2 U648 ( .A(\r524/A[0] ), .B(\eq_112/B[0] ), .Z(n864) );
  NOR4_X2 U649 ( .A1(n868), .A2(n869), .A3(n870), .A4(n871), .ZN(n862) );
  XOR2_X2 U650 ( .A(\r524/A[7] ), .B(\eq_112/B[7] ), .Z(n871) );
  XOR2_X2 U651 ( .A(\r524/A[6] ), .B(\eq_112/B[6] ), .Z(n870) );
  XOR2_X2 U652 ( .A(\r524/A[5] ), .B(\eq_112/B[5] ), .Z(n869) );
  XOR2_X2 U653 ( .A(\r524/A[4] ), .B(\eq_112/B[4] ), .Z(n868) );
  NOR4_X2 U654 ( .A1(n872), .A2(n873), .A3(n874), .A4(n875), .ZN(n861) );
  XOR2_X2 U655 ( .A(\r524/A[11] ), .B(\eq_112/B[11] ), .Z(n875) );
  XOR2_X2 U656 ( .A(\r524/A[10] ), .B(\eq_112/B[10] ), .Z(n874) );
  XOR2_X2 U657 ( .A(\r524/A[9] ), .B(\eq_112/B[9] ), .Z(n873) );
  XOR2_X2 U658 ( .A(\r524/A[8] ), .B(\eq_112/B[8] ), .Z(n872) );
  NOR4_X2 U659 ( .A1(n876), .A2(n877), .A3(n878), .A4(n879), .ZN(n860) );
  XOR2_X2 U660 ( .A(\r524/A[15] ), .B(\eq_112/B[15] ), .Z(n879) );
  XOR2_X2 U661 ( .A(\r524/A[14] ), .B(\eq_112/B[14] ), .Z(n878) );
  XOR2_X2 U662 ( .A(\r524/A[13] ), .B(\eq_112/B[13] ), .Z(n877) );
  XOR2_X2 U663 ( .A(\r524/A[12] ), .B(\eq_112/B[12] ), .Z(n876) );
  NAND4_X2 U664 ( .A1(n880), .A2(n881), .A3(n882), .A4(n883), .ZN(n822) );
  NOR4_X2 U665 ( .A1(n884), .A2(n885), .A3(n886), .A4(n887), .ZN(n883) );
  XOR2_X2 U666 ( .A(\r523/A[3] ), .B(\eq_112/B[3] ), .Z(n887) );
  XOR2_X2 U667 ( .A(\r523/A[2] ), .B(\eq_112/B[2] ), .Z(n886) );
  XOR2_X2 U668 ( .A(\r523/A[1] ), .B(\eq_112/B[1] ), .Z(n885) );
  XOR2_X2 U669 ( .A(\r523/A[0] ), .B(\eq_112/B[0] ), .Z(n884) );
  NOR4_X2 U670 ( .A1(n888), .A2(n889), .A3(n890), .A4(n891), .ZN(n882) );
  XOR2_X2 U671 ( .A(\r523/A[7] ), .B(\eq_112/B[7] ), .Z(n891) );
  XOR2_X2 U672 ( .A(\r523/A[6] ), .B(\eq_112/B[6] ), .Z(n890) );
  XOR2_X2 U673 ( .A(\r523/A[5] ), .B(\eq_112/B[5] ), .Z(n889) );
  XOR2_X2 U674 ( .A(\r523/A[4] ), .B(\eq_112/B[4] ), .Z(n888) );
  NOR4_X2 U675 ( .A1(n892), .A2(n893), .A3(n894), .A4(n895), .ZN(n881) );
  XOR2_X2 U676 ( .A(\r523/A[11] ), .B(\eq_112/B[11] ), .Z(n895) );
  XOR2_X2 U677 ( .A(\r523/A[10] ), .B(\eq_112/B[10] ), .Z(n894) );
  XOR2_X2 U678 ( .A(\r523/A[9] ), .B(\eq_112/B[9] ), .Z(n893) );
  XOR2_X2 U679 ( .A(\r523/A[8] ), .B(\eq_112/B[8] ), .Z(n892) );
  NOR4_X2 U680 ( .A1(n896), .A2(n897), .A3(n898), .A4(n899), .ZN(n880) );
  XOR2_X2 U681 ( .A(\r523/A[15] ), .B(\eq_112/B[15] ), .Z(n899) );
  XOR2_X2 U682 ( .A(\r523/A[14] ), .B(\eq_112/B[14] ), .Z(n898) );
  XOR2_X2 U683 ( .A(\r523/A[13] ), .B(\eq_112/B[13] ), .Z(n897) );
  XOR2_X2 U684 ( .A(\r523/A[12] ), .B(\eq_112/B[12] ), .Z(n896) );
  NAND4_X2 U685 ( .A1(n900), .A2(n901), .A3(n902), .A4(n903), .ZN(n821) );
  NOR4_X2 U686 ( .A1(n904), .A2(n905), .A3(n906), .A4(n907), .ZN(n903) );
  XOR2_X2 U687 ( .A(\eq_112/B[3] ), .B(\eq_112/A[3] ), .Z(n907) );
  XOR2_X2 U688 ( .A(\eq_112/B[2] ), .B(\eq_112/A[2] ), .Z(n906) );
  XOR2_X2 U689 ( .A(\eq_112/B[1] ), .B(\eq_112/A[1] ), .Z(n905) );
  XOR2_X2 U690 ( .A(\eq_112/B[0] ), .B(\eq_112/A[0] ), .Z(n904) );
  NOR4_X2 U691 ( .A1(n908), .A2(n909), .A3(n910), .A4(n911), .ZN(n902) );
  XOR2_X2 U692 ( .A(\eq_112/B[7] ), .B(\eq_112/A[7] ), .Z(n911) );
  XOR2_X2 U693 ( .A(\eq_112/B[6] ), .B(\eq_112/A[6] ), .Z(n910) );
  XOR2_X2 U694 ( .A(\eq_112/B[5] ), .B(\eq_112/A[5] ), .Z(n909) );
  XOR2_X2 U695 ( .A(\eq_112/B[4] ), .B(\eq_112/A[4] ), .Z(n908) );
  NOR4_X2 U696 ( .A1(n912), .A2(n913), .A3(n914), .A4(n915), .ZN(n901) );
  XOR2_X2 U697 ( .A(\eq_112/B[11] ), .B(\eq_112/A[11] ), .Z(n915) );
  XOR2_X2 U698 ( .A(\eq_112/B[10] ), .B(\eq_112/A[10] ), .Z(n914) );
  XOR2_X2 U699 ( .A(\eq_112/B[9] ), .B(\eq_112/A[9] ), .Z(n913) );
  XOR2_X2 U700 ( .A(\eq_112/B[8] ), .B(\eq_112/A[8] ), .Z(n912) );
  NOR4_X2 U701 ( .A1(n916), .A2(n917), .A3(n918), .A4(n919), .ZN(n900) );
  XOR2_X2 U702 ( .A(\eq_112/B[15] ), .B(\eq_112/A[15] ), .Z(n919) );
  XOR2_X2 U703 ( .A(\eq_112/B[14] ), .B(\eq_112/A[14] ), .Z(n918) );
  XOR2_X2 U704 ( .A(\eq_112/B[13] ), .B(\eq_112/A[13] ), .Z(n917) );
  XOR2_X2 U705 ( .A(\eq_112/B[12] ), .B(\eq_112/A[12] ), .Z(n916) );
  NAND2_X2 U707 ( .A1(PosRowY[1]), .A2(n921), .ZN(n922) );
  OAI221_X2 U710 ( .B1(n3962), .B2(n3939), .C1(n834), .C2(n925), .A(n212), 
        .ZN(n924) );
  NAND2_X2 U711 ( .A1(n3963), .A2(n3939), .ZN(n212) );
  NAND2_X2 U712 ( .A1(n925), .A2(n926), .ZN(n833) );
  NAND2_X2 U726 ( .A1(n825), .A2(n3919), .ZN(n831) );
  OAI22_X2 U727 ( .A1(n29), .A2(n938), .B1(n3957), .B2(n3921), .ZN(n1078) );
  NAND3_X2 U729 ( .A1(n3963), .A2(n3958), .A3(PosDY[1]), .ZN(n940) );
  NOR2_X2 U731 ( .A1(n3958), .A2(PosDY[1]), .ZN(n805) );
  NOR2_X2 U732 ( .A1(PosDY[1]), .A2(PosDY[0]), .ZN(n807) );
  NAND2_X2 U733 ( .A1(n832), .A2(n825), .ZN(n938) );
  NAND3_X2 U735 ( .A1(DiagonalDoneY), .A2(n28), .A3(FoundY[0]), .ZN(n827) );
  NAND2_X2 U736 ( .A1(n920), .A2(n834), .ZN(n823) );
  NAND4_X2 U737 ( .A1(n943), .A2(n944), .A3(n945), .A4(n946), .ZN(n834) );
  NOR4_X2 U738 ( .A1(n947), .A2(n948), .A3(n949), .A4(n950), .ZN(n946) );
  XOR2_X2 U739 ( .A(\r526/A[3] ), .B(\eq_207/B[3] ), .Z(n950) );
  XOR2_X2 U740 ( .A(\r526/A[2] ), .B(\eq_207/B[2] ), .Z(n949) );
  XOR2_X2 U741 ( .A(\r526/A[1] ), .B(\eq_207/B[1] ), .Z(n948) );
  XOR2_X2 U742 ( .A(\r526/A[0] ), .B(\eq_207/B[0] ), .Z(n947) );
  NOR4_X2 U743 ( .A1(n951), .A2(n952), .A3(n953), .A4(n954), .ZN(n945) );
  XOR2_X2 U744 ( .A(\r526/A[7] ), .B(\eq_207/B[7] ), .Z(n954) );
  XOR2_X2 U745 ( .A(\r526/A[6] ), .B(\eq_207/B[6] ), .Z(n953) );
  XOR2_X2 U746 ( .A(\r526/A[5] ), .B(\eq_207/B[5] ), .Z(n952) );
  XOR2_X2 U747 ( .A(\r526/A[4] ), .B(\eq_207/B[4] ), .Z(n951) );
  NOR4_X2 U748 ( .A1(n955), .A2(n956), .A3(n957), .A4(n958), .ZN(n944) );
  XOR2_X2 U749 ( .A(\r526/A[11] ), .B(\eq_207/B[11] ), .Z(n958) );
  XOR2_X2 U750 ( .A(\r526/A[10] ), .B(\eq_207/B[10] ), .Z(n957) );
  XOR2_X2 U751 ( .A(\r526/A[9] ), .B(\eq_207/B[9] ), .Z(n956) );
  XOR2_X2 U752 ( .A(\r526/A[8] ), .B(\eq_207/B[8] ), .Z(n955) );
  NOR4_X2 U753 ( .A1(n959), .A2(n960), .A3(n961), .A4(n962), .ZN(n943) );
  XOR2_X2 U754 ( .A(\r526/A[15] ), .B(\eq_207/B[15] ), .Z(n962) );
  XOR2_X2 U755 ( .A(\r526/A[14] ), .B(\eq_207/B[14] ), .Z(n961) );
  XOR2_X2 U756 ( .A(\r526/A[13] ), .B(\eq_207/B[13] ), .Z(n960) );
  XOR2_X2 U757 ( .A(\r526/A[12] ), .B(\eq_207/B[12] ), .Z(n959) );
  NOR2_X2 U758 ( .A1(n925), .A2(n3963), .ZN(n920) );
  NAND4_X2 U759 ( .A1(n963), .A2(n964), .A3(n965), .A4(n966), .ZN(n926) );
  NOR4_X2 U760 ( .A1(n967), .A2(n968), .A3(n969), .A4(n970), .ZN(n966) );
  XOR2_X2 U761 ( .A(\r528/A[3] ), .B(\eq_207/B[3] ), .Z(n970) );
  XOR2_X2 U762 ( .A(\r528/A[2] ), .B(\eq_207/B[2] ), .Z(n969) );
  XOR2_X2 U763 ( .A(\r528/A[1] ), .B(\eq_207/B[1] ), .Z(n968) );
  XOR2_X2 U764 ( .A(\r528/A[0] ), .B(\eq_207/B[0] ), .Z(n967) );
  NOR4_X2 U765 ( .A1(n971), .A2(n972), .A3(n973), .A4(n974), .ZN(n965) );
  XOR2_X2 U766 ( .A(\r528/A[7] ), .B(\eq_207/B[7] ), .Z(n974) );
  XOR2_X2 U767 ( .A(\r528/A[6] ), .B(\eq_207/B[6] ), .Z(n973) );
  XOR2_X2 U768 ( .A(\r528/A[5] ), .B(\eq_207/B[5] ), .Z(n972) );
  XOR2_X2 U769 ( .A(\r528/A[4] ), .B(\eq_207/B[4] ), .Z(n971) );
  NOR4_X2 U770 ( .A1(n975), .A2(n976), .A3(n977), .A4(n978), .ZN(n964) );
  XOR2_X2 U771 ( .A(\r528/A[11] ), .B(\eq_207/B[11] ), .Z(n978) );
  XOR2_X2 U772 ( .A(\r528/A[10] ), .B(\eq_207/B[10] ), .Z(n977) );
  XOR2_X2 U773 ( .A(\r528/A[9] ), .B(\eq_207/B[9] ), .Z(n976) );
  XOR2_X2 U774 ( .A(\r528/A[8] ), .B(\eq_207/B[8] ), .Z(n975) );
  NOR4_X2 U775 ( .A1(n979), .A2(n980), .A3(n981), .A4(n982), .ZN(n963) );
  XOR2_X2 U776 ( .A(\r528/A[15] ), .B(\eq_207/B[15] ), .Z(n982) );
  XOR2_X2 U777 ( .A(\r528/A[14] ), .B(\eq_207/B[14] ), .Z(n981) );
  XOR2_X2 U778 ( .A(\r528/A[13] ), .B(\eq_207/B[13] ), .Z(n980) );
  XOR2_X2 U779 ( .A(\r528/A[12] ), .B(\eq_207/B[12] ), .Z(n979) );
  AND4_X2 U780 ( .A1(n983), .A2(n984), .A3(n985), .A4(n986), .ZN(n925) );
  NOR4_X2 U781 ( .A1(n987), .A2(n988), .A3(n989), .A4(n990), .ZN(n986) );
  XOR2_X2 U782 ( .A(\r527/A[3] ), .B(\eq_207/B[3] ), .Z(n990) );
  XOR2_X2 U783 ( .A(\r527/A[2] ), .B(\eq_207/B[2] ), .Z(n989) );
  XOR2_X2 U784 ( .A(\r527/A[1] ), .B(\eq_207/B[1] ), .Z(n988) );
  XOR2_X2 U785 ( .A(\r527/A[0] ), .B(\eq_207/B[0] ), .Z(n987) );
  NOR4_X2 U786 ( .A1(n991), .A2(n992), .A3(n993), .A4(n994), .ZN(n985) );
  XOR2_X2 U787 ( .A(\r527/A[7] ), .B(\eq_207/B[7] ), .Z(n994) );
  XOR2_X2 U788 ( .A(\r527/A[6] ), .B(\eq_207/B[6] ), .Z(n993) );
  XOR2_X2 U789 ( .A(\r527/A[5] ), .B(\eq_207/B[5] ), .Z(n992) );
  XOR2_X2 U790 ( .A(\r527/A[4] ), .B(\eq_207/B[4] ), .Z(n991) );
  NOR4_X2 U791 ( .A1(n995), .A2(n996), .A3(n997), .A4(n998), .ZN(n984) );
  XOR2_X2 U792 ( .A(\r527/A[11] ), .B(\eq_207/B[11] ), .Z(n998) );
  XOR2_X2 U793 ( .A(\r527/A[10] ), .B(\eq_207/B[10] ), .Z(n997) );
  XOR2_X2 U794 ( .A(\r527/A[9] ), .B(\eq_207/B[9] ), .Z(n996) );
  XOR2_X2 U795 ( .A(\r527/A[8] ), .B(\eq_207/B[8] ), .Z(n995) );
  NOR4_X2 U796 ( .A1(n999), .A2(n1000), .A3(n1001), .A4(n1002), .ZN(n983) );
  XOR2_X2 U797 ( .A(\r527/A[15] ), .B(\eq_207/B[15] ), .Z(n1002) );
  XOR2_X2 U798 ( .A(\r527/A[14] ), .B(\eq_207/B[14] ), .Z(n1001) );
  XOR2_X2 U799 ( .A(\r527/A[13] ), .B(\eq_207/B[13] ), .Z(n1000) );
  XOR2_X2 U800 ( .A(\r527/A[12] ), .B(\eq_207/B[12] ), .Z(n999) );
  NAND4_X2 U801 ( .A1(n1003), .A2(n1004), .A3(n1005), .A4(n1006), .ZN(n826) );
  NOR4_X2 U802 ( .A1(n1007), .A2(n1008), .A3(n1009), .A4(n1010), .ZN(n1006) );
  XOR2_X2 U803 ( .A(\eq_207/B[3] ), .B(\eq_207/A[3] ), .Z(n1010) );
  XOR2_X2 U804 ( .A(\eq_207/B[2] ), .B(\eq_207/A[2] ), .Z(n1009) );
  XOR2_X2 U805 ( .A(\eq_207/B[1] ), .B(\eq_207/A[1] ), .Z(n1008) );
  XOR2_X2 U806 ( .A(\eq_207/B[0] ), .B(\eq_207/A[0] ), .Z(n1007) );
  NOR4_X2 U807 ( .A1(n1011), .A2(n1012), .A3(n1013), .A4(n1014), .ZN(n1005) );
  XOR2_X2 U808 ( .A(\eq_207/B[7] ), .B(\eq_207/A[7] ), .Z(n1014) );
  XOR2_X2 U809 ( .A(\eq_207/B[6] ), .B(\eq_207/A[6] ), .Z(n1013) );
  XOR2_X2 U810 ( .A(\eq_207/B[5] ), .B(\eq_207/A[5] ), .Z(n1012) );
  XOR2_X2 U811 ( .A(\eq_207/B[4] ), .B(\eq_207/A[4] ), .Z(n1011) );
  NOR4_X2 U812 ( .A1(n1015), .A2(n1016), .A3(n1017), .A4(n1018), .ZN(n1004) );
  XOR2_X2 U813 ( .A(\eq_207/B[11] ), .B(\eq_207/A[11] ), .Z(n1018) );
  XOR2_X2 U814 ( .A(\eq_207/B[10] ), .B(\eq_207/A[10] ), .Z(n1017) );
  XOR2_X2 U815 ( .A(\eq_207/B[9] ), .B(\eq_207/A[9] ), .Z(n1016) );
  XOR2_X2 U816 ( .A(\eq_207/B[8] ), .B(\eq_207/A[8] ), .Z(n1015) );
  NOR4_X2 U817 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1003) );
  XOR2_X2 U818 ( .A(\eq_207/B[15] ), .B(\eq_207/A[15] ), .Z(n1022) );
  XOR2_X2 U819 ( .A(\eq_207/B[14] ), .B(\eq_207/A[14] ), .Z(n1021) );
  XOR2_X2 U820 ( .A(\eq_207/B[13] ), .B(\eq_207/A[13] ), .Z(n1020) );
  XOR2_X2 U821 ( .A(\eq_207/B[12] ), .B(\eq_207/A[12] ), .Z(n1019) );
  NOR2_X2 U822 ( .A1(reset), .A2(EnableChange), .ZN(n832) );
  NAND3_X2 U824 ( .A1(n29), .A2(n28), .A3(DiagonalDoneY), .ZN(n939) );
  NAND3_X2 U826 ( .A1(n36), .A2(n35), .A3(DiagonalDoneX), .ZN(n836) );
  AND2_X1 U1015 ( .A1(n231), .A2(n232), .ZN(n221) );
  AND2_X1 U1016 ( .A1(n254), .A2(n255), .ZN(n251) );
  AND2_X1 U1017 ( .A1(n266), .A2(n267), .ZN(n263) );
  AND2_X1 U1018 ( .A1(n278), .A2(n279), .ZN(n275) );
  AND2_X1 U1019 ( .A1(n290), .A2(n291), .ZN(n287) );
  AND2_X1 U1020 ( .A1(n302), .A2(n303), .ZN(n299) );
  AND2_X1 U1021 ( .A1(n314), .A2(n315), .ZN(n311) );
  AND2_X1 U1022 ( .A1(n326), .A2(n327), .ZN(n323) );
  AND2_X1 U1023 ( .A1(n338), .A2(n339), .ZN(n335) );
  AND2_X1 U1024 ( .A1(n350), .A2(n351), .ZN(n347) );
  AND2_X1 U1025 ( .A1(n362), .A2(n363), .ZN(n359) );
  AND2_X1 U1026 ( .A1(n374), .A2(n375), .ZN(n371) );
  AND2_X1 U1027 ( .A1(n386), .A2(n387), .ZN(n383) );
  AND2_X1 U1028 ( .A1(n398), .A2(n399), .ZN(n395) );
  AND2_X1 U1029 ( .A1(n410), .A2(n411), .ZN(n407) );
  AND2_X1 U1030 ( .A1(n422), .A2(n423), .ZN(n419) );
  AND2_X1 U1031 ( .A1(n434), .A2(n435), .ZN(n431) );
  AND2_X1 U1032 ( .A1(n446), .A2(n447), .ZN(n443) );
  AND2_X1 U1033 ( .A1(n458), .A2(n459), .ZN(n455) );
  AND2_X1 U1034 ( .A1(n470), .A2(n471), .ZN(n467) );
  AND2_X1 U1035 ( .A1(n482), .A2(n483), .ZN(n479) );
  AND2_X1 U1036 ( .A1(n494), .A2(n495), .ZN(n491) );
  AND2_X1 U1037 ( .A1(n506), .A2(n507), .ZN(n503) );
  AND2_X1 U1038 ( .A1(n518), .A2(n519), .ZN(n515) );
  AND2_X1 U1039 ( .A1(n530), .A2(n531), .ZN(n527) );
  AND2_X1 U1040 ( .A1(n542), .A2(n543), .ZN(n539) );
  AND2_X1 U1041 ( .A1(n554), .A2(n555), .ZN(n551) );
  AND2_X1 U1042 ( .A1(n566), .A2(n567), .ZN(n563) );
  AND2_X1 U1043 ( .A1(n578), .A2(n579), .ZN(n575) );
  AND2_X1 U1044 ( .A1(n590), .A2(n591), .ZN(n587) );
  AND2_X1 U1045 ( .A1(n602), .A2(n603), .ZN(n599) );
  AND2_X1 U1046 ( .A1(n614), .A2(n615), .ZN(n611) );
  AND2_X1 U1047 ( .A1(n626), .A2(n627), .ZN(n623) );
  AND2_X1 U1048 ( .A1(n638), .A2(n639), .ZN(n635) );
  AND2_X1 U1049 ( .A1(n650), .A2(n651), .ZN(n647) );
  AND2_X1 U1050 ( .A1(n662), .A2(n663), .ZN(n659) );
  AND2_X1 U1051 ( .A1(n674), .A2(n675), .ZN(n671) );
  AND2_X1 U1052 ( .A1(n686), .A2(n687), .ZN(n683) );
  AND2_X1 U1053 ( .A1(n698), .A2(n699), .ZN(n695) );
  AND2_X1 U1054 ( .A1(n710), .A2(n711), .ZN(n707) );
  AND2_X1 U1055 ( .A1(n722), .A2(n723), .ZN(n719) );
  AND2_X1 U1056 ( .A1(n734), .A2(n735), .ZN(n731) );
  AND2_X1 U1057 ( .A1(n746), .A2(n747), .ZN(n743) );
  AND2_X1 U1058 ( .A1(n758), .A2(n759), .ZN(n755) );
  AND2_X1 U1059 ( .A1(n770), .A2(n771), .ZN(n767) );
  AND2_X1 U1060 ( .A1(n782), .A2(n783), .ZN(n779) );
  AND2_X1 U1061 ( .A1(n794), .A2(n795), .ZN(n791) );
  AND2_X1 U1066 ( .A1(n809), .A2(n810), .ZN(n803) );
  AND2_X1 U1076 ( .A1(n3965), .A2(n817), .ZN(n839) );
  OR2_X1 U1077 ( .A1(n939), .A2(n940), .ZN(n220) );
  AND2_X1 U1078 ( .A1(n3961), .A2(n805), .ZN(n942) );
  DFF_X2 \FoundY_reg[1]  ( .D(n1077), .CK(clock), .Q(FoundY[1]), .QN(n28) );
  DFF_X2 \FoundX_reg[1]  ( .D(n1073), .CK(clock), .Q(FoundX[1]), .QN(n35) );
  OR2_X4 U3 ( .A1(n926), .A2(n827), .ZN(n3924) );
  OR2_X4 U5 ( .A1(n939), .A2(n940), .ZN(n3919) );
  MUX2_X2 U6 ( .A(PosRowX[0]), .B(n196), .S(n201), .Z(n1024) );
  MUX2_X2 U8 ( .A(n924), .B(PosRowY[0]), .S(n921), .Z(n1076) );
  AND2_X4 U9 ( .A1(n824), .A2(n825), .ZN(n3889) );
  AND2_X4 U10 ( .A1(n805), .A2(n3962), .ZN(n3890) );
  AND2_X4 U11 ( .A1(n805), .A2(n3963), .ZN(n3891) );
  AND2_X4 U12 ( .A1(n807), .A2(n808), .ZN(n3892) );
  AND2_X4 U13 ( .A1(n807), .A2(n823), .ZN(n3893) );
  AND2_X4 U14 ( .A1(n197), .A2(n3954), .ZN(n3894) );
  NOR2_X4 U15 ( .A1(n833), .A2(n827), .ZN(n3895) );
  OR2_X4 U16 ( .A1(n836), .A2(n838), .ZN(n3896) );
  NAND2_X4 U17 ( .A1(n817), .A2(n813), .ZN(n3897) );
  AND2_X4 U18 ( .A1(n816), .A2(n815), .ZN(n3898) );
  NAND2_X4 U19 ( .A1(n197), .A2(n817), .ZN(n3899) );
  AND2_X4 U20 ( .A1(n815), .A2(n813), .ZN(n3900) );
  NOR3_X4 U21 ( .A1(n819), .A2(n820), .A3(n821), .ZN(n3901) );
  AND2_X4 U22 ( .A1(n807), .A2(n3962), .ZN(n3902) );
  AND2_X4 U24 ( .A1(n197), .A2(n815), .ZN(n242) );
  AND2_X4 U26 ( .A1(WireY), .A2(n940), .ZN(n3903) );
  NAND2_X2 U28 ( .A1(n816), .A2(n3954), .ZN(n3904) );
  AND2_X4 U29 ( .A1(n3954), .A2(n813), .ZN(n3905) );
  NAND2_X2 U30 ( .A1(n3939), .A2(n808), .ZN(n3906) );
  INV_X4 U31 ( .A(n3905), .ZN(n3926) );
  INV_X4 U32 ( .A(n818), .ZN(n3910) );
  INV_X4 U33 ( .A(n3904), .ZN(n3913) );
  INV_X4 U34 ( .A(n3904), .ZN(n3914) );
  INV_X4 U36 ( .A(n3906), .ZN(n3911) );
  INV_X4 U38 ( .A(n3906), .ZN(n3912) );
  INV_X4 U40 ( .A(n3905), .ZN(n3925) );
  INV_X4 U41 ( .A(n3923), .ZN(n3922) );
  INV_X4 U42 ( .A(n3903), .ZN(n3920) );
  INV_X4 U43 ( .A(n3903), .ZN(n3921) );
  INV_X4 U44 ( .A(n3915), .ZN(n3916) );
  INV_X4 U45 ( .A(n939), .ZN(WireY) );
  OAI21_X2 U46 ( .B1(n3964), .B2(n820), .A(n3954), .ZN(n828) );
  OAI21_X2 U48 ( .B1(n3960), .B2(n823), .A(n3939), .ZN(n825) );
  INV_X4 U50 ( .A(n215), .ZN(n3923) );
  INV_X4 U52 ( .A(n921), .ZN(n3907) );
  AOI21_X2 U53 ( .B1(WireY), .B2(n3957), .A(n831), .ZN(n921) );
  INV_X4 U54 ( .A(n201), .ZN(n3953) );
  INV_X4 U55 ( .A(n3918), .ZN(n3917) );
  INV_X4 U56 ( .A(n222), .ZN(n3918) );
  INV_X4 U57 ( .A(n939), .ZN(n3908) );
  AOI222_X1 U58 ( .A1(n804), .A2(n222), .B1(\U93/DATA1_0 ), .B2(n3890), .C1(
        \U90/DATA1_0 ), .C2(n3891), .ZN(n802) );
  AOI22_X2 U60 ( .A1(\U95/DATA1_0 ), .A2(n3892), .B1(\U93/DATA1_0 ), .B2(n3902), .ZN(n806) );
  AOI222_X1 U62 ( .A1(n792), .A2(n222), .B1(\U93/DATA1_1 ), .B2(n3890), .C1(
        \U90/DATA1_1 ), .C2(n3891), .ZN(n790) );
  AOI22_X2 U64 ( .A1(\U95/DATA1_1 ), .A2(n3892), .B1(\U93/DATA1_1 ), .B2(n3902), .ZN(n793) );
  AOI222_X1 U65 ( .A1(n780), .A2(n3917), .B1(\U93/DATA1_2 ), .B2(n3890), .C1(
        \U90/DATA1_2 ), .C2(n3891), .ZN(n778) );
  AOI22_X2 U66 ( .A1(\U95/DATA1_2 ), .A2(n3892), .B1(\U93/DATA1_2 ), .B2(n3902), .ZN(n781) );
  AOI222_X1 U67 ( .A1(n768), .A2(n222), .B1(\U93/DATA1_3 ), .B2(n3890), .C1(
        \U90/DATA1_3 ), .C2(n3891), .ZN(n766) );
  AOI22_X2 U68 ( .A1(\U95/DATA1_3 ), .A2(n3892), .B1(\U93/DATA1_3 ), .B2(n3902), .ZN(n769) );
  AOI222_X1 U69 ( .A1(n756), .A2(n222), .B1(\U93/DATA1_4 ), .B2(n3890), .C1(
        \U90/DATA1_4 ), .C2(n3891), .ZN(n754) );
  AOI22_X2 U70 ( .A1(\U95/DATA1_4 ), .A2(n3892), .B1(\U93/DATA1_4 ), .B2(n3902), .ZN(n757) );
  AOI222_X1 U72 ( .A1(n744), .A2(n3917), .B1(\U93/DATA1_5 ), .B2(n3890), .C1(
        \U90/DATA1_5 ), .C2(n3891), .ZN(n742) );
  AOI22_X2 U74 ( .A1(\U95/DATA1_5 ), .A2(n3892), .B1(\U93/DATA1_5 ), .B2(n3902), .ZN(n745) );
  AOI222_X1 U76 ( .A1(n732), .A2(n222), .B1(\U93/DATA1_6 ), .B2(n3890), .C1(
        \U90/DATA1_6 ), .C2(n3891), .ZN(n730) );
  AOI22_X2 U77 ( .A1(\U95/DATA1_6 ), .A2(n3892), .B1(\U93/DATA1_6 ), .B2(n3902), .ZN(n733) );
  AOI222_X1 U78 ( .A1(n720), .A2(n222), .B1(\U93/DATA1_7 ), .B2(n3890), .C1(
        \U90/DATA1_7 ), .C2(n3891), .ZN(n718) );
  AOI22_X2 U79 ( .A1(\U95/DATA1_7 ), .A2(n3892), .B1(\U93/DATA1_7 ), .B2(n3902), .ZN(n721) );
  AOI222_X1 U80 ( .A1(n708), .A2(n222), .B1(\U93/DATA1_8 ), .B2(n3890), .C1(
        \U90/DATA1_8 ), .C2(n3891), .ZN(n706) );
  AOI22_X2 U81 ( .A1(\U95/DATA1_8 ), .A2(n3892), .B1(\U93/DATA1_8 ), .B2(n3902), .ZN(n709) );
  AOI222_X1 U82 ( .A1(n696), .A2(n3917), .B1(\U93/DATA1_9 ), .B2(n3890), .C1(
        \U90/DATA1_9 ), .C2(n3891), .ZN(n694) );
  AOI22_X2 U84 ( .A1(\U95/DATA1_9 ), .A2(n3892), .B1(\U93/DATA1_9 ), .B2(n3902), .ZN(n697) );
  AOI222_X1 U86 ( .A1(n684), .A2(n3917), .B1(\U93/DATA1_10 ), .B2(n3890), .C1(
        \U90/DATA1_10 ), .C2(n3891), .ZN(n682) );
  AOI22_X2 U88 ( .A1(\U95/DATA1_10 ), .A2(n3892), .B1(\U93/DATA1_10 ), .B2(
        n3902), .ZN(n685) );
  AOI222_X1 U89 ( .A1(n672), .A2(n3917), .B1(\U93/DATA1_11 ), .B2(n3890), .C1(
        \U90/DATA1_11 ), .C2(n3891), .ZN(n670) );
  AOI22_X2 U90 ( .A1(\U95/DATA1_11 ), .A2(n3892), .B1(\U93/DATA1_11 ), .B2(
        n3902), .ZN(n673) );
  AOI222_X1 U91 ( .A1(n648), .A2(n3917), .B1(\U93/DATA1_13 ), .B2(n3890), .C1(
        \U90/DATA1_13 ), .C2(n3891), .ZN(n646) );
  AOI22_X2 U92 ( .A1(\U95/DATA1_13 ), .A2(n3892), .B1(\U93/DATA1_13 ), .B2(
        n3902), .ZN(n649) );
  AOI222_X1 U93 ( .A1(n636), .A2(n222), .B1(\U93/DATA1_14 ), .B2(n3890), .C1(
        \U90/DATA1_14 ), .C2(n3891), .ZN(n634) );
  AOI22_X2 U94 ( .A1(\U95/DATA1_14 ), .A2(n3892), .B1(\U93/DATA1_14 ), .B2(
        n3902), .ZN(n637) );
  AOI222_X1 U96 ( .A1(n624), .A2(n222), .B1(\U93/DATA1_15 ), .B2(n3890), .C1(
        \U90/DATA1_15 ), .C2(n3891), .ZN(n622) );
  AOI22_X2 U98 ( .A1(\U95/DATA1_15 ), .A2(n3892), .B1(\U93/DATA1_15 ), .B2(
        n3902), .ZN(n625) );
  AOI222_X1 U100 ( .A1(n612), .A2(n222), .B1(\U93/DATA1_16 ), .B2(n3890), .C1(
        \U90/DATA1_16 ), .C2(n3891), .ZN(n610) );
  AOI22_X2 U101 ( .A1(\U95/DATA1_16 ), .A2(n3892), .B1(\U93/DATA1_16 ), .B2(
        n3902), .ZN(n613) );
  AOI222_X1 U102 ( .A1(n600), .A2(n222), .B1(\U93/DATA1_17 ), .B2(n3890), .C1(
        \U90/DATA1_17 ), .C2(n3891), .ZN(n598) );
  AOI22_X2 U103 ( .A1(\U95/DATA1_17 ), .A2(n3892), .B1(\U93/DATA1_17 ), .B2(
        n3902), .ZN(n601) );
  AOI222_X1 U104 ( .A1(n588), .A2(n222), .B1(\U93/DATA1_18 ), .B2(n3890), .C1(
        \U90/DATA1_18 ), .C2(n3891), .ZN(n586) );
  AOI22_X2 U105 ( .A1(\U95/DATA1_18 ), .A2(n3892), .B1(\U93/DATA1_18 ), .B2(
        n3902), .ZN(n589) );
  AOI222_X1 U106 ( .A1(n576), .A2(n222), .B1(\U93/DATA1_19 ), .B2(n3890), .C1(
        \U90/DATA1_19 ), .C2(n3891), .ZN(n574) );
  AOI22_X2 U108 ( .A1(\U95/DATA1_19 ), .A2(n3892), .B1(\U93/DATA1_19 ), .B2(
        n3902), .ZN(n577) );
  AOI222_X1 U110 ( .A1(n564), .A2(n222), .B1(\U93/DATA1_20 ), .B2(n3890), .C1(
        \U90/DATA1_20 ), .C2(n3891), .ZN(n562) );
  AOI22_X2 U112 ( .A1(\U95/DATA1_20 ), .A2(n3892), .B1(\U93/DATA1_20 ), .B2(
        n3902), .ZN(n565) );
  AOI222_X1 U113 ( .A1(n552), .A2(n222), .B1(\U93/DATA1_21 ), .B2(n3890), .C1(
        \U90/DATA1_21 ), .C2(n3891), .ZN(n550) );
  AOI22_X2 U114 ( .A1(\U95/DATA1_21 ), .A2(n3892), .B1(\U93/DATA1_21 ), .B2(
        n3902), .ZN(n553) );
  AOI222_X1 U115 ( .A1(n540), .A2(n222), .B1(\U93/DATA1_22 ), .B2(n3890), .C1(
        \U90/DATA1_22 ), .C2(n3891), .ZN(n538) );
  AOI22_X2 U116 ( .A1(\U95/DATA1_22 ), .A2(n3892), .B1(\U93/DATA1_22 ), .B2(
        n3902), .ZN(n541) );
  AOI222_X1 U117 ( .A1(n528), .A2(n222), .B1(\U93/DATA1_23 ), .B2(n3890), .C1(
        \U90/DATA1_23 ), .C2(n3891), .ZN(n526) );
  AOI22_X2 U118 ( .A1(\U95/DATA1_23 ), .A2(n3892), .B1(\U93/DATA1_23 ), .B2(
        n3902), .ZN(n529) );
  AOI222_X1 U120 ( .A1(n516), .A2(n222), .B1(\U93/DATA1_24 ), .B2(n3890), .C1(
        \U90/DATA1_24 ), .C2(n3891), .ZN(n514) );
  AOI22_X2 U122 ( .A1(\U95/DATA1_24 ), .A2(n3892), .B1(\U93/DATA1_24 ), .B2(
        n3902), .ZN(n517) );
  AOI222_X1 U124 ( .A1(n504), .A2(n222), .B1(\U93/DATA1_25 ), .B2(n3890), .C1(
        \U90/DATA1_25 ), .C2(n3891), .ZN(n502) );
  AOI22_X2 U125 ( .A1(\U95/DATA1_25 ), .A2(n3892), .B1(\U93/DATA1_25 ), .B2(
        n3902), .ZN(n505) );
  AOI222_X1 U126 ( .A1(n492), .A2(n222), .B1(\U93/DATA1_26 ), .B2(n3890), .C1(
        \U90/DATA1_26 ), .C2(n3891), .ZN(n490) );
  AOI22_X2 U127 ( .A1(\U95/DATA1_26 ), .A2(n3892), .B1(\U93/DATA1_26 ), .B2(
        n3902), .ZN(n493) );
  AOI222_X1 U128 ( .A1(n480), .A2(n222), .B1(\U93/DATA1_27 ), .B2(n3890), .C1(
        \U90/DATA1_27 ), .C2(n3891), .ZN(n478) );
  AOI22_X2 U129 ( .A1(\U95/DATA1_27 ), .A2(n3892), .B1(\U93/DATA1_27 ), .B2(
        n3902), .ZN(n481) );
  AOI222_X1 U130 ( .A1(n468), .A2(n222), .B1(\U93/DATA1_28 ), .B2(n3890), .C1(
        \U90/DATA1_28 ), .C2(n3891), .ZN(n466) );
  AOI22_X2 U132 ( .A1(\U95/DATA1_28 ), .A2(n3892), .B1(\U93/DATA1_28 ), .B2(
        n3902), .ZN(n469) );
  AOI222_X1 U134 ( .A1(n456), .A2(n222), .B1(\U93/DATA1_29 ), .B2(n3890), .C1(
        \U90/DATA1_29 ), .C2(n3891), .ZN(n454) );
  AOI22_X2 U136 ( .A1(\U95/DATA1_29 ), .A2(n3892), .B1(\U93/DATA1_29 ), .B2(
        n3902), .ZN(n457) );
  AOI222_X1 U137 ( .A1(n444), .A2(n222), .B1(\U93/DATA1_30 ), .B2(n3890), .C1(
        \U90/DATA1_30 ), .C2(n3891), .ZN(n442) );
  AOI22_X2 U138 ( .A1(\U95/DATA1_30 ), .A2(n3892), .B1(\U93/DATA1_30 ), .B2(
        n3902), .ZN(n445) );
  AOI222_X1 U139 ( .A1(n432), .A2(n222), .B1(\U93/DATA1_31 ), .B2(n3890), .C1(
        \U90/DATA1_31 ), .C2(n3891), .ZN(n430) );
  AOI22_X2 U140 ( .A1(\U95/DATA1_31 ), .A2(n3892), .B1(\U93/DATA1_31 ), .B2(
        n3902), .ZN(n433) );
  AOI222_X1 U141 ( .A1(n420), .A2(n222), .B1(\U93/DATA1_32 ), .B2(n3890), .C1(
        \U90/DATA1_32 ), .C2(n3891), .ZN(n418) );
  AOI22_X2 U142 ( .A1(\U95/DATA1_32 ), .A2(n3892), .B1(\U93/DATA1_32 ), .B2(
        n3902), .ZN(n421) );
  AOI222_X1 U144 ( .A1(n408), .A2(n222), .B1(\U93/DATA1_33 ), .B2(n3890), .C1(
        \U90/DATA1_33 ), .C2(n3891), .ZN(n406) );
  AOI22_X2 U146 ( .A1(\U95/DATA1_33 ), .A2(n3892), .B1(\U93/DATA1_33 ), .B2(
        n3902), .ZN(n409) );
  AOI222_X1 U148 ( .A1(n396), .A2(n222), .B1(\U93/DATA1_34 ), .B2(n3890), .C1(
        \U90/DATA1_34 ), .C2(n3891), .ZN(n394) );
  AOI22_X2 U149 ( .A1(\U95/DATA1_34 ), .A2(n3892), .B1(\U93/DATA1_34 ), .B2(
        n3902), .ZN(n397) );
  AOI222_X1 U150 ( .A1(n384), .A2(n3917), .B1(\U93/DATA1_35 ), .B2(n3890), 
        .C1(\U90/DATA1_35 ), .C2(n3891), .ZN(n382) );
  AOI22_X2 U151 ( .A1(\U95/DATA1_35 ), .A2(n3892), .B1(\U93/DATA1_35 ), .B2(
        n3902), .ZN(n385) );
  AOI222_X1 U152 ( .A1(n372), .A2(n3917), .B1(\U93/DATA1_36 ), .B2(n3890), 
        .C1(\U90/DATA1_36 ), .C2(n3891), .ZN(n370) );
  AOI22_X2 U153 ( .A1(\U95/DATA1_36 ), .A2(n3892), .B1(\U93/DATA1_36 ), .B2(
        n3902), .ZN(n373) );
  AOI222_X1 U154 ( .A1(n360), .A2(n3917), .B1(\U93/DATA1_37 ), .B2(n3890), 
        .C1(\U90/DATA1_37 ), .C2(n3891), .ZN(n358) );
  AOI22_X2 U156 ( .A1(\U95/DATA1_37 ), .A2(n3892), .B1(\U93/DATA1_37 ), .B2(
        n3902), .ZN(n361) );
  AOI222_X1 U158 ( .A1(n348), .A2(n3917), .B1(\U93/DATA1_38 ), .B2(n3890), 
        .C1(\U90/DATA1_38 ), .C2(n3891), .ZN(n346) );
  AOI22_X2 U160 ( .A1(\U95/DATA1_38 ), .A2(n3892), .B1(\U93/DATA1_38 ), .B2(
        n3902), .ZN(n349) );
  AOI222_X1 U161 ( .A1(n336), .A2(n3917), .B1(\U93/DATA1_39 ), .B2(n3890), 
        .C1(\U90/DATA1_39 ), .C2(n3891), .ZN(n334) );
  AOI22_X2 U162 ( .A1(\U95/DATA1_39 ), .A2(n3892), .B1(\U93/DATA1_39 ), .B2(
        n3902), .ZN(n337) );
  AOI222_X1 U163 ( .A1(n324), .A2(n3917), .B1(\U93/DATA1_40 ), .B2(n3890), 
        .C1(\U90/DATA1_40 ), .C2(n3891), .ZN(n322) );
  AOI22_X2 U164 ( .A1(\U95/DATA1_40 ), .A2(n3892), .B1(\U93/DATA1_40 ), .B2(
        n3902), .ZN(n325) );
  AOI222_X1 U165 ( .A1(n312), .A2(n3917), .B1(\U93/DATA1_41 ), .B2(n3890), 
        .C1(\U90/DATA1_41 ), .C2(n3891), .ZN(n310) );
  AOI22_X2 U166 ( .A1(\U95/DATA1_41 ), .A2(n3892), .B1(\U93/DATA1_41 ), .B2(
        n3902), .ZN(n313) );
  AOI222_X1 U168 ( .A1(n300), .A2(n3917), .B1(\U93/DATA1_42 ), .B2(n3890), 
        .C1(\U90/DATA1_42 ), .C2(n3891), .ZN(n298) );
  AOI22_X2 U170 ( .A1(\U95/DATA1_42 ), .A2(n3892), .B1(\U93/DATA1_42 ), .B2(
        n3902), .ZN(n301) );
  AOI222_X1 U172 ( .A1(n288), .A2(n3917), .B1(\U93/DATA1_43 ), .B2(n3890), 
        .C1(\U90/DATA1_43 ), .C2(n3891), .ZN(n286) );
  AOI22_X2 U173 ( .A1(\U95/DATA1_43 ), .A2(n3892), .B1(\U93/DATA1_43 ), .B2(
        n3902), .ZN(n289) );
  AOI222_X1 U174 ( .A1(n276), .A2(n3917), .B1(\U93/DATA1_44 ), .B2(n3890), 
        .C1(\U90/DATA1_44 ), .C2(n3891), .ZN(n274) );
  AOI22_X2 U175 ( .A1(\U95/DATA1_44 ), .A2(n3892), .B1(\U93/DATA1_44 ), .B2(
        n3902), .ZN(n277) );
  AOI222_X1 U176 ( .A1(n264), .A2(n3917), .B1(\U93/DATA1_45 ), .B2(n3890), 
        .C1(\U90/DATA1_45 ), .C2(n3891), .ZN(n262) );
  AOI22_X2 U177 ( .A1(\U95/DATA1_45 ), .A2(n3892), .B1(\U93/DATA1_45 ), .B2(
        n3902), .ZN(n265) );
  AOI222_X1 U178 ( .A1(n252), .A2(n3917), .B1(\U93/DATA1_46 ), .B2(n3890), 
        .C1(\U90/DATA1_46 ), .C2(n3891), .ZN(n250) );
  AOI22_X2 U180 ( .A1(\U95/DATA1_46 ), .A2(n3892), .B1(\U93/DATA1_46 ), .B2(
        n3902), .ZN(n253) );
  AOI222_X1 U182 ( .A1(n660), .A2(n222), .B1(\U93/DATA1_12 ), .B2(n3890), .C1(
        \U90/DATA1_12 ), .C2(n3891), .ZN(n658) );
  AOI22_X2 U184 ( .A1(\U95/DATA1_12 ), .A2(n3892), .B1(\U93/DATA1_12 ), .B2(
        n3902), .ZN(n661) );
  AOI222_X1 U185 ( .A1(n3917), .A2(n223), .B1(n3890), .B2(\U93/DATA1_47 ), 
        .C1(n3891), .C2(\U90/DATA1_47 ), .ZN(n218) );
  AOI22_X2 U186 ( .A1(n3892), .A2(\U95/DATA1_47 ), .B1(n3902), .B2(
        \U93/DATA1_47 ), .ZN(n228) );
  AOI222_X1 U187 ( .A1(\U163/DATA1_0 ), .A2(n3900), .B1(\U168/DATA1_0 ), .B2(
        n3898), .C1(\U166/DATA1_0 ), .C2(n242), .ZN(n814) );
  AOI222_X1 U188 ( .A1(\U163/DATA1_1 ), .A2(n3900), .B1(\U168/DATA1_1 ), .B2(
        n3898), .C1(\U166/DATA1_1 ), .C2(n242), .ZN(n798) );
  AOI222_X1 U189 ( .A1(\U163/DATA1_2 ), .A2(n3900), .B1(\U168/DATA1_2 ), .B2(
        n3898), .C1(\U166/DATA1_2 ), .C2(n242), .ZN(n786) );
  AOI222_X1 U190 ( .A1(\U163/DATA1_3 ), .A2(n3900), .B1(\U168/DATA1_3 ), .B2(
        n3898), .C1(\U166/DATA1_3 ), .C2(n242), .ZN(n774) );
  AOI222_X1 U192 ( .A1(\U163/DATA1_4 ), .A2(n3900), .B1(\U168/DATA1_4 ), .B2(
        n3898), .C1(\U166/DATA1_4 ), .C2(n242), .ZN(n762) );
  AOI222_X1 U194 ( .A1(\U163/DATA1_5 ), .A2(n3900), .B1(\U168/DATA1_5 ), .B2(
        n3898), .C1(\U166/DATA1_5 ), .C2(n242), .ZN(n750) );
  AOI222_X1 U196 ( .A1(\U163/DATA1_6 ), .A2(n3900), .B1(\U168/DATA1_6 ), .B2(
        n3898), .C1(\U166/DATA1_6 ), .C2(n242), .ZN(n738) );
  AOI222_X1 U197 ( .A1(\U163/DATA1_7 ), .A2(n3900), .B1(\U168/DATA1_7 ), .B2(
        n3898), .C1(\U166/DATA1_7 ), .C2(n242), .ZN(n726) );
  AOI222_X1 U198 ( .A1(\U163/DATA1_8 ), .A2(n3900), .B1(\U168/DATA1_8 ), .B2(
        n3898), .C1(\U166/DATA1_8 ), .C2(n242), .ZN(n714) );
  AOI222_X1 U199 ( .A1(\U163/DATA1_9 ), .A2(n3900), .B1(\U168/DATA1_9 ), .B2(
        n3898), .C1(\U166/DATA1_9 ), .C2(n242), .ZN(n702) );
  AOI222_X1 U200 ( .A1(\U163/DATA1_10 ), .A2(n3900), .B1(\U168/DATA1_10 ), 
        .B2(n3898), .C1(\U166/DATA1_10 ), .C2(n242), .ZN(n690) );
  AOI222_X1 U201 ( .A1(\U163/DATA1_11 ), .A2(n3900), .B1(\U168/DATA1_11 ), 
        .B2(n3898), .C1(\U166/DATA1_11 ), .C2(n242), .ZN(n678) );
  AOI222_X1 U202 ( .A1(\U163/DATA1_12 ), .A2(n3900), .B1(\U168/DATA1_12 ), 
        .B2(n3898), .C1(\U166/DATA1_12 ), .C2(n242), .ZN(n666) );
  AOI222_X1 U204 ( .A1(\U163/DATA1_13 ), .A2(n3900), .B1(\U168/DATA1_13 ), 
        .B2(n3898), .C1(\U166/DATA1_13 ), .C2(n242), .ZN(n654) );
  AOI222_X1 U206 ( .A1(\U163/DATA1_14 ), .A2(n3900), .B1(\U168/DATA1_14 ), 
        .B2(n3898), .C1(\U166/DATA1_14 ), .C2(n242), .ZN(n642) );
  AOI222_X1 U208 ( .A1(\U163/DATA1_15 ), .A2(n3900), .B1(\U168/DATA1_15 ), 
        .B2(n3898), .C1(\U166/DATA1_15 ), .C2(n242), .ZN(n630) );
  AOI222_X1 U209 ( .A1(\U163/DATA1_16 ), .A2(n3900), .B1(\U168/DATA1_16 ), 
        .B2(n3898), .C1(\U166/DATA1_16 ), .C2(n242), .ZN(n618) );
  AOI222_X1 U210 ( .A1(\U163/DATA1_17 ), .A2(n3900), .B1(\U168/DATA1_17 ), 
        .B2(n3898), .C1(\U166/DATA1_17 ), .C2(n242), .ZN(n606) );
  AOI222_X1 U211 ( .A1(\U163/DATA1_18 ), .A2(n3900), .B1(\U168/DATA1_18 ), 
        .B2(n3898), .C1(\U166/DATA1_18 ), .C2(n242), .ZN(n594) );
  AOI222_X1 U212 ( .A1(\U163/DATA1_19 ), .A2(n3900), .B1(\U168/DATA1_19 ), 
        .B2(n3898), .C1(\U166/DATA1_19 ), .C2(n242), .ZN(n582) );
  AOI222_X1 U213 ( .A1(\U163/DATA1_20 ), .A2(n3900), .B1(\U168/DATA1_20 ), 
        .B2(n3898), .C1(\U166/DATA1_20 ), .C2(n242), .ZN(n570) );
  AOI222_X1 U214 ( .A1(\U163/DATA1_21 ), .A2(n3900), .B1(\U168/DATA1_21 ), 
        .B2(n3898), .C1(\U166/DATA1_21 ), .C2(n242), .ZN(n558) );
  AOI222_X1 U216 ( .A1(\U163/DATA1_22 ), .A2(n3900), .B1(\U168/DATA1_22 ), 
        .B2(n3898), .C1(\U166/DATA1_22 ), .C2(n242), .ZN(n546) );
  AOI222_X1 U218 ( .A1(\U163/DATA1_23 ), .A2(n3900), .B1(\U168/DATA1_23 ), 
        .B2(n3898), .C1(\U166/DATA1_23 ), .C2(n242), .ZN(n534) );
  AOI222_X1 U220 ( .A1(\U163/DATA1_24 ), .A2(n3900), .B1(\U168/DATA1_24 ), 
        .B2(n3898), .C1(\U166/DATA1_24 ), .C2(n242), .ZN(n522) );
  AOI222_X1 U221 ( .A1(\U163/DATA1_25 ), .A2(n3900), .B1(\U168/DATA1_25 ), 
        .B2(n3898), .C1(\U166/DATA1_25 ), .C2(n242), .ZN(n510) );
  AOI222_X1 U222 ( .A1(\U163/DATA1_26 ), .A2(n3900), .B1(\U168/DATA1_26 ), 
        .B2(n3898), .C1(\U166/DATA1_26 ), .C2(n242), .ZN(n498) );
  AOI222_X1 U223 ( .A1(\U163/DATA1_27 ), .A2(n3900), .B1(\U168/DATA1_27 ), 
        .B2(n3898), .C1(\U166/DATA1_27 ), .C2(n242), .ZN(n486) );
  AOI222_X1 U224 ( .A1(\U163/DATA1_28 ), .A2(n3900), .B1(\U168/DATA1_28 ), 
        .B2(n3898), .C1(\U166/DATA1_28 ), .C2(n242), .ZN(n474) );
  AOI222_X1 U225 ( .A1(\U163/DATA1_29 ), .A2(n3900), .B1(\U168/DATA1_29 ), 
        .B2(n3898), .C1(\U166/DATA1_29 ), .C2(n242), .ZN(n462) );
  AOI222_X1 U226 ( .A1(\U163/DATA1_30 ), .A2(n3900), .B1(\U168/DATA1_30 ), 
        .B2(n3898), .C1(\U166/DATA1_30 ), .C2(n242), .ZN(n450) );
  AOI222_X1 U228 ( .A1(\U163/DATA1_31 ), .A2(n3900), .B1(\U168/DATA1_31 ), 
        .B2(n3898), .C1(\U166/DATA1_31 ), .C2(n242), .ZN(n438) );
  AOI222_X1 U230 ( .A1(\U163/DATA1_32 ), .A2(n3900), .B1(\U168/DATA1_32 ), 
        .B2(n3898), .C1(\U166/DATA1_32 ), .C2(n242), .ZN(n426) );
  AOI222_X1 U232 ( .A1(\U163/DATA1_33 ), .A2(n3900), .B1(\U168/DATA1_33 ), 
        .B2(n3898), .C1(\U166/DATA1_33 ), .C2(n242), .ZN(n414) );
  AOI222_X1 U233 ( .A1(\U163/DATA1_34 ), .A2(n3900), .B1(\U168/DATA1_34 ), 
        .B2(n3898), .C1(\U166/DATA1_34 ), .C2(n242), .ZN(n402) );
  AOI222_X1 U234 ( .A1(\U163/DATA1_47 ), .A2(n3900), .B1(\U168/DATA1_47 ), 
        .B2(n3898), .C1(\U166/DATA1_47 ), .C2(n242), .ZN(n239) );
  AOI222_X1 U235 ( .A1(\U163/DATA1_35 ), .A2(n3900), .B1(\U168/DATA1_35 ), 
        .B2(n3898), .C1(\U166/DATA1_35 ), .C2(n242), .ZN(n390) );
  AOI222_X1 U236 ( .A1(\U163/DATA1_36 ), .A2(n3900), .B1(\U168/DATA1_36 ), 
        .B2(n3898), .C1(\U166/DATA1_36 ), .C2(n242), .ZN(n378) );
  AOI222_X1 U237 ( .A1(\U163/DATA1_37 ), .A2(n3900), .B1(\U168/DATA1_37 ), 
        .B2(n3898), .C1(\U166/DATA1_37 ), .C2(n242), .ZN(n366) );
  AOI222_X1 U238 ( .A1(\U163/DATA1_38 ), .A2(n3900), .B1(\U168/DATA1_38 ), 
        .B2(n3898), .C1(\U166/DATA1_38 ), .C2(n242), .ZN(n354) );
  AOI222_X1 U240 ( .A1(\U163/DATA1_39 ), .A2(n3900), .B1(\U168/DATA1_39 ), 
        .B2(n3898), .C1(\U166/DATA1_39 ), .C2(n242), .ZN(n342) );
  AOI222_X1 U242 ( .A1(\U163/DATA1_40 ), .A2(n3900), .B1(\U168/DATA1_40 ), 
        .B2(n3898), .C1(\U166/DATA1_40 ), .C2(n242), .ZN(n330) );
  AOI222_X1 U244 ( .A1(\U163/DATA1_41 ), .A2(n3900), .B1(\U168/DATA1_41 ), 
        .B2(n3898), .C1(\U166/DATA1_41 ), .C2(n242), .ZN(n318) );
  AOI222_X1 U245 ( .A1(\U163/DATA1_42 ), .A2(n3900), .B1(\U168/DATA1_42 ), 
        .B2(n3898), .C1(\U166/DATA1_42 ), .C2(n242), .ZN(n306) );
  AOI222_X1 U246 ( .A1(\U163/DATA1_43 ), .A2(n3900), .B1(\U168/DATA1_43 ), 
        .B2(n3898), .C1(\U166/DATA1_43 ), .C2(n242), .ZN(n294) );
  AOI222_X1 U247 ( .A1(\U163/DATA1_44 ), .A2(n3900), .B1(\U168/DATA1_44 ), 
        .B2(n3898), .C1(\U166/DATA1_44 ), .C2(n242), .ZN(n282) );
  AOI222_X1 U248 ( .A1(\U163/DATA1_45 ), .A2(n3900), .B1(\U168/DATA1_45 ), 
        .B2(n3898), .C1(\U166/DATA1_45 ), .C2(n242), .ZN(n270) );
  AOI222_X1 U249 ( .A1(\U163/DATA1_46 ), .A2(n3900), .B1(\U168/DATA1_46 ), 
        .B2(n3898), .C1(\U166/DATA1_46 ), .C2(n242), .ZN(n258) );
  AOI22_X2 U250 ( .A1(n3894), .A2(\U166/DATA1_47 ), .B1(\U125/DATA1_47 ), .B2(
        n3901), .ZN(n231) );
  AOI21_X2 U252 ( .B1(n3925), .B2(n3896), .A(n4015), .ZN(n235) );
  AOI22_X2 U254 ( .A1(\U166/DATA1_0 ), .A2(n3894), .B1(\U125/DATA1_0 ), .B2(
        n3901), .ZN(n809) );
  AOI21_X2 U256 ( .B1(n3925), .B2(n3896), .A(n4062), .ZN(n812) );
  AOI22_X2 U257 ( .A1(\U166/DATA1_1 ), .A2(n3894), .B1(\U125/DATA1_1 ), .B2(
        n3901), .ZN(n794) );
  AOI21_X2 U258 ( .B1(n3925), .B2(n3896), .A(n4061), .ZN(n797) );
  AOI22_X2 U259 ( .A1(\U166/DATA1_2 ), .A2(n3894), .B1(\U125/DATA1_2 ), .B2(
        n3901), .ZN(n782) );
  AOI21_X2 U260 ( .B1(n3925), .B2(n3896), .A(n4060), .ZN(n785) );
  AOI22_X2 U261 ( .A1(\U166/DATA1_3 ), .A2(n3894), .B1(\U125/DATA1_3 ), .B2(
        n3901), .ZN(n770) );
  AOI21_X2 U262 ( .B1(n3925), .B2(n3896), .A(n4059), .ZN(n773) );
  AOI22_X2 U264 ( .A1(\U166/DATA1_4 ), .A2(n3894), .B1(\U125/DATA1_4 ), .B2(
        n3901), .ZN(n758) );
  AOI21_X2 U266 ( .B1(n3925), .B2(n3896), .A(n4058), .ZN(n761) );
  AOI22_X2 U268 ( .A1(\U166/DATA1_5 ), .A2(n3894), .B1(\U125/DATA1_5 ), .B2(
        n3901), .ZN(n746) );
  AOI21_X2 U269 ( .B1(n3925), .B2(n3896), .A(n4057), .ZN(n749) );
  AOI22_X2 U270 ( .A1(\U166/DATA1_6 ), .A2(n3894), .B1(\U125/DATA1_6 ), .B2(
        n3901), .ZN(n734) );
  AOI21_X2 U271 ( .B1(n3925), .B2(n3896), .A(n4056), .ZN(n737) );
  AOI22_X2 U272 ( .A1(\U166/DATA1_7 ), .A2(n3894), .B1(\U125/DATA1_7 ), .B2(
        n3901), .ZN(n722) );
  AOI21_X2 U273 ( .B1(n3925), .B2(n3896), .A(n4055), .ZN(n725) );
  AOI22_X2 U274 ( .A1(\U166/DATA1_8 ), .A2(n3894), .B1(\U125/DATA1_8 ), .B2(
        n3901), .ZN(n710) );
  AOI21_X2 U276 ( .B1(n3925), .B2(n3896), .A(n4054), .ZN(n713) );
  AOI22_X2 U278 ( .A1(\U166/DATA1_9 ), .A2(n3894), .B1(\U125/DATA1_9 ), .B2(
        n3901), .ZN(n698) );
  AOI21_X2 U280 ( .B1(n3925), .B2(n3896), .A(n4053), .ZN(n701) );
  AOI22_X2 U281 ( .A1(\U166/DATA1_10 ), .A2(n3894), .B1(\U125/DATA1_10 ), .B2(
        n3901), .ZN(n686) );
  AOI21_X2 U282 ( .B1(n3925), .B2(n3896), .A(n4052), .ZN(n689) );
  AOI22_X2 U283 ( .A1(\U166/DATA1_11 ), .A2(n3894), .B1(\U125/DATA1_11 ), .B2(
        n3901), .ZN(n674) );
  AOI21_X2 U284 ( .B1(n3925), .B2(n3896), .A(n4051), .ZN(n677) );
  AOI22_X2 U285 ( .A1(\U166/DATA1_12 ), .A2(n3894), .B1(\U125/DATA1_12 ), .B2(
        n3901), .ZN(n662) );
  AOI21_X2 U286 ( .B1(n3925), .B2(n3896), .A(n4050), .ZN(n665) );
  AOI22_X2 U288 ( .A1(\U166/DATA1_13 ), .A2(n3894), .B1(\U125/DATA1_13 ), .B2(
        n3901), .ZN(n650) );
  AOI21_X2 U290 ( .B1(n3926), .B2(n3896), .A(n4049), .ZN(n653) );
  AOI22_X2 U292 ( .A1(\U166/DATA1_14 ), .A2(n3894), .B1(\U125/DATA1_14 ), .B2(
        n3901), .ZN(n638) );
  AOI21_X2 U293 ( .B1(n3926), .B2(n3896), .A(n4048), .ZN(n641) );
  AOI22_X2 U294 ( .A1(\U166/DATA1_15 ), .A2(n3894), .B1(\U125/DATA1_15 ), .B2(
        n3901), .ZN(n626) );
  AOI21_X2 U295 ( .B1(n3926), .B2(n3896), .A(n4047), .ZN(n629) );
  AOI22_X2 U296 ( .A1(\U166/DATA1_16 ), .A2(n3894), .B1(\U125/DATA1_16 ), .B2(
        n3901), .ZN(n614) );
  AOI21_X2 U297 ( .B1(n3926), .B2(n3896), .A(n4046), .ZN(n617) );
  AOI22_X2 U298 ( .A1(\U166/DATA1_17 ), .A2(n3894), .B1(\U125/DATA1_17 ), .B2(
        n3901), .ZN(n602) );
  AOI21_X2 U300 ( .B1(n3926), .B2(n3896), .A(n4045), .ZN(n605) );
  AOI22_X2 U302 ( .A1(\U166/DATA1_18 ), .A2(n3894), .B1(\U125/DATA1_18 ), .B2(
        n3901), .ZN(n590) );
  AOI21_X2 U304 ( .B1(n3925), .B2(n3896), .A(n4044), .ZN(n593) );
  AOI22_X2 U305 ( .A1(\U166/DATA1_19 ), .A2(n3894), .B1(\U125/DATA1_19 ), .B2(
        n3901), .ZN(n578) );
  AOI21_X2 U306 ( .B1(n3926), .B2(n3896), .A(n4043), .ZN(n581) );
  AOI22_X2 U307 ( .A1(\U166/DATA1_20 ), .A2(n3894), .B1(\U125/DATA1_20 ), .B2(
        n3901), .ZN(n566) );
  AOI21_X2 U308 ( .B1(n3925), .B2(n3896), .A(n4042), .ZN(n569) );
  AOI22_X2 U309 ( .A1(\U166/DATA1_21 ), .A2(n3894), .B1(\U125/DATA1_21 ), .B2(
        n3901), .ZN(n554) );
  AOI21_X2 U310 ( .B1(n3926), .B2(n3896), .A(n4041), .ZN(n557) );
  AOI22_X2 U312 ( .A1(\U166/DATA1_22 ), .A2(n3894), .B1(\U125/DATA1_22 ), .B2(
        n3901), .ZN(n542) );
  AOI21_X2 U314 ( .B1(n3925), .B2(n3896), .A(n4040), .ZN(n545) );
  AOI22_X2 U316 ( .A1(\U166/DATA1_23 ), .A2(n3894), .B1(\U125/DATA1_23 ), .B2(
        n3901), .ZN(n530) );
  AOI21_X2 U317 ( .B1(n3926), .B2(n3896), .A(n4039), .ZN(n533) );
  AOI22_X2 U318 ( .A1(\U166/DATA1_24 ), .A2(n3894), .B1(\U125/DATA1_24 ), .B2(
        n3901), .ZN(n518) );
  AOI21_X2 U319 ( .B1(n3925), .B2(n3896), .A(n4038), .ZN(n521) );
  AOI22_X2 U320 ( .A1(\U166/DATA1_25 ), .A2(n3894), .B1(\U125/DATA1_25 ), .B2(
        n3901), .ZN(n506) );
  AOI21_X2 U321 ( .B1(n3926), .B2(n3896), .A(n4037), .ZN(n509) );
  AOI22_X2 U322 ( .A1(\U166/DATA1_26 ), .A2(n3894), .B1(\U125/DATA1_26 ), .B2(
        n3901), .ZN(n494) );
  AOI21_X2 U324 ( .B1(n3926), .B2(n3896), .A(n4036), .ZN(n497) );
  AOI22_X2 U326 ( .A1(\U166/DATA1_27 ), .A2(n3894), .B1(\U125/DATA1_27 ), .B2(
        n3901), .ZN(n482) );
  AOI21_X2 U328 ( .B1(n3926), .B2(n3896), .A(n4035), .ZN(n485) );
  AOI22_X2 U329 ( .A1(\U166/DATA1_28 ), .A2(n3894), .B1(\U125/DATA1_28 ), .B2(
        n3901), .ZN(n470) );
  AOI21_X2 U330 ( .B1(n3926), .B2(n3896), .A(n4034), .ZN(n473) );
  AOI22_X2 U331 ( .A1(\U166/DATA1_29 ), .A2(n3894), .B1(\U125/DATA1_29 ), .B2(
        n3901), .ZN(n458) );
  AOI21_X2 U332 ( .B1(n3926), .B2(n3896), .A(n4033), .ZN(n461) );
  AOI22_X2 U333 ( .A1(\U166/DATA1_30 ), .A2(n3894), .B1(\U125/DATA1_30 ), .B2(
        n3901), .ZN(n446) );
  AOI21_X2 U334 ( .B1(n3926), .B2(n3896), .A(n4032), .ZN(n449) );
  AOI22_X2 U336 ( .A1(\U166/DATA1_31 ), .A2(n3894), .B1(\U125/DATA1_31 ), .B2(
        n3901), .ZN(n434) );
  AOI21_X2 U338 ( .B1(n3926), .B2(n3896), .A(n4031), .ZN(n437) );
  AOI22_X2 U340 ( .A1(\U166/DATA1_32 ), .A2(n3894), .B1(\U125/DATA1_32 ), .B2(
        n3901), .ZN(n422) );
  AOI21_X2 U341 ( .B1(n3926), .B2(n3896), .A(n4030), .ZN(n425) );
  AOI22_X2 U342 ( .A1(\U166/DATA1_33 ), .A2(n3894), .B1(\U125/DATA1_33 ), .B2(
        n3901), .ZN(n410) );
  AOI21_X2 U343 ( .B1(n3926), .B2(n3896), .A(n4029), .ZN(n413) );
  AOI22_X2 U344 ( .A1(\U166/DATA1_34 ), .A2(n3894), .B1(\U125/DATA1_34 ), .B2(
        n3901), .ZN(n398) );
  AOI21_X2 U345 ( .B1(n3926), .B2(n3896), .A(n4028), .ZN(n401) );
  AOI22_X2 U346 ( .A1(\U166/DATA1_35 ), .A2(n3894), .B1(\U125/DATA1_35 ), .B2(
        n3901), .ZN(n386) );
  AOI21_X2 U348 ( .B1(n3926), .B2(n3896), .A(n4027), .ZN(n389) );
  AOI22_X2 U350 ( .A1(\U166/DATA1_36 ), .A2(n3894), .B1(\U125/DATA1_36 ), .B2(
        n3901), .ZN(n374) );
  AOI21_X2 U352 ( .B1(n3926), .B2(n3896), .A(n4026), .ZN(n377) );
  AOI22_X2 U353 ( .A1(\U166/DATA1_37 ), .A2(n3894), .B1(\U125/DATA1_37 ), .B2(
        n3901), .ZN(n362) );
  AOI21_X2 U354 ( .B1(n3926), .B2(n3896), .A(n4025), .ZN(n365) );
  AOI22_X2 U355 ( .A1(\U166/DATA1_38 ), .A2(n3894), .B1(\U125/DATA1_38 ), .B2(
        n3901), .ZN(n350) );
  AOI21_X2 U356 ( .B1(n3926), .B2(n3896), .A(n4024), .ZN(n353) );
  AOI22_X2 U357 ( .A1(\U166/DATA1_39 ), .A2(n3894), .B1(\U125/DATA1_39 ), .B2(
        n3901), .ZN(n338) );
  AOI21_X2 U358 ( .B1(n3926), .B2(n3896), .A(n4023), .ZN(n341) );
  AOI22_X2 U360 ( .A1(\U166/DATA1_40 ), .A2(n3894), .B1(\U125/DATA1_40 ), .B2(
        n3901), .ZN(n326) );
  AOI21_X2 U362 ( .B1(n3925), .B2(n3896), .A(n4022), .ZN(n329) );
  AOI22_X2 U364 ( .A1(\U166/DATA1_41 ), .A2(n3894), .B1(\U125/DATA1_41 ), .B2(
        n3901), .ZN(n314) );
  AOI21_X2 U365 ( .B1(n3926), .B2(n3896), .A(n4021), .ZN(n317) );
  AOI22_X2 U366 ( .A1(\U166/DATA1_42 ), .A2(n3894), .B1(\U125/DATA1_42 ), .B2(
        n3901), .ZN(n302) );
  AOI21_X2 U367 ( .B1(n3925), .B2(n3896), .A(n4020), .ZN(n305) );
  AOI22_X2 U368 ( .A1(\U166/DATA1_43 ), .A2(n3894), .B1(\U125/DATA1_43 ), .B2(
        n3901), .ZN(n290) );
  AOI21_X2 U369 ( .B1(n3926), .B2(n3896), .A(n4019), .ZN(n293) );
  AOI22_X2 U370 ( .A1(\U166/DATA1_44 ), .A2(n3894), .B1(\U125/DATA1_44 ), .B2(
        n3901), .ZN(n278) );
  AOI21_X2 U372 ( .B1(n3925), .B2(n3896), .A(n4018), .ZN(n281) );
  AOI22_X2 U374 ( .A1(\U166/DATA1_45 ), .A2(n3894), .B1(\U125/DATA1_45 ), .B2(
        n3901), .ZN(n266) );
  AOI21_X2 U376 ( .B1(n3926), .B2(n3896), .A(n4017), .ZN(n269) );
  AOI22_X2 U377 ( .A1(\U166/DATA1_46 ), .A2(n3894), .B1(\U125/DATA1_46 ), .B2(
        n3901), .ZN(n254) );
  AOI21_X2 U378 ( .B1(n3925), .B2(n3896), .A(n4016), .ZN(n257) );
  AOI211_X2 U379 ( .C1(n3957), .C2(n3908), .A(n831), .B(n3959), .ZN(n830) );
  OAI21_X2 U380 ( .B1(n815), .B2(n839), .A(n820), .ZN(n837) );
  OAI21_X2 U381 ( .B1(n807), .B2(n942), .A(n823), .ZN(n941) );
  OAI211_X2 U382 ( .C1(n836), .C2(n837), .A(n828), .B(n3896), .ZN(n201) );
  INV_X4 U384 ( .A(n226), .ZN(n3915) );
  OAI211_X2 U386 ( .C1(n3924), .C2(n4098), .A(n655), .B(n656), .ZN(n1060) );
  AOI22_X2 U388 ( .A1(\U95/DATA1_12 ), .A2(n3911), .B1(\U93/DATA1_12 ), .B2(
        n3895), .ZN(n655) );
  AOI222_X1 U389 ( .A1(Element[12]), .A2(n3927), .B1(\U52/DATA1_12 ), .B2(
        n3922), .C1(n3889), .C2(n657), .ZN(n656) );
  OAI222_X2 U390 ( .A1(n658), .A2(n3921), .B1(n220), .B2(n4098), .C1(WireY), 
        .C2(n659), .ZN(n657) );
  OAI211_X2 U391 ( .C1(n3924), .C2(n4097), .A(n643), .B(n644), .ZN(n1059) );
  AOI22_X2 U392 ( .A1(\U95/DATA1_13 ), .A2(n3911), .B1(\U93/DATA1_13 ), .B2(
        n3895), .ZN(n643) );
  AOI222_X1 U393 ( .A1(Element[13]), .A2(n3927), .B1(\U52/DATA1_13 ), .B2(
        n3922), .C1(n3889), .C2(n645), .ZN(n644) );
  OAI222_X2 U394 ( .A1(n646), .A2(n3920), .B1(n220), .B2(n4097), .C1(WireY), 
        .C2(n647), .ZN(n645) );
  OAI211_X2 U396 ( .C1(n3924), .C2(n4096), .A(n631), .B(n632), .ZN(n1058) );
  AOI22_X2 U398 ( .A1(\U95/DATA1_14 ), .A2(n3911), .B1(\U93/DATA1_14 ), .B2(
        n3895), .ZN(n631) );
  AOI222_X1 U400 ( .A1(Element[14]), .A2(n3927), .B1(\U52/DATA1_14 ), .B2(
        n3922), .C1(n3889), .C2(n633), .ZN(n632) );
  OAI222_X2 U401 ( .A1(n634), .A2(n3921), .B1(n220), .B2(n4096), .C1(WireY), 
        .C2(n635), .ZN(n633) );
  OAI211_X2 U402 ( .C1(n3924), .C2(n4095), .A(n619), .B(n620), .ZN(n1057) );
  AOI22_X2 U403 ( .A1(\U95/DATA1_15 ), .A2(n3911), .B1(\U93/DATA1_15 ), .B2(
        n3895), .ZN(n619) );
  AOI222_X1 U404 ( .A1(Element[15]), .A2(n3927), .B1(\U52/DATA1_15 ), .B2(
        n3922), .C1(n3889), .C2(n621), .ZN(n620) );
  OAI222_X2 U405 ( .A1(n622), .A2(n3920), .B1(n220), .B2(n4095), .C1(WireY), 
        .C2(n623), .ZN(n621) );
  OAI211_X2 U406 ( .C1(n3924), .C2(n4094), .A(n607), .B(n608), .ZN(n1056) );
  AOI22_X2 U408 ( .A1(\U95/DATA1_16 ), .A2(n3911), .B1(\U93/DATA1_16 ), .B2(
        n3895), .ZN(n607) );
  AOI222_X1 U410 ( .A1(Element[16]), .A2(n3927), .B1(\U52/DATA1_16 ), .B2(
        n3922), .C1(n3889), .C2(n609), .ZN(n608) );
  OAI222_X2 U412 ( .A1(n610), .A2(n3921), .B1(n220), .B2(n4094), .C1(WireY), 
        .C2(n611), .ZN(n609) );
  OAI211_X2 U413 ( .C1(n3924), .C2(n4093), .A(n595), .B(n596), .ZN(n1055) );
  AOI22_X2 U414 ( .A1(\U95/DATA1_17 ), .A2(n3911), .B1(\U93/DATA1_17 ), .B2(
        n3895), .ZN(n595) );
  AOI222_X1 U415 ( .A1(Element[17]), .A2(n3927), .B1(\U52/DATA1_17 ), .B2(
        n3922), .C1(n3889), .C2(n597), .ZN(n596) );
  OAI222_X2 U416 ( .A1(n598), .A2(n3920), .B1(n220), .B2(n4093), .C1(WireY), 
        .C2(n599), .ZN(n597) );
  OAI211_X2 U417 ( .C1(n3924), .C2(n4092), .A(n583), .B(n584), .ZN(n1054) );
  AOI22_X2 U418 ( .A1(\U95/DATA1_18 ), .A2(n3911), .B1(\U93/DATA1_18 ), .B2(
        n3895), .ZN(n583) );
  AOI222_X1 U420 ( .A1(Element[18]), .A2(n3927), .B1(\U52/DATA1_18 ), .B2(
        n3922), .C1(n3889), .C2(n585), .ZN(n584) );
  OAI222_X2 U422 ( .A1(n586), .A2(n3921), .B1(n220), .B2(n4092), .C1(WireY), 
        .C2(n587), .ZN(n585) );
  OAI211_X2 U424 ( .C1(n3924), .C2(n4091), .A(n571), .B(n572), .ZN(n1053) );
  AOI22_X2 U425 ( .A1(\U95/DATA1_19 ), .A2(n3911), .B1(\U93/DATA1_19 ), .B2(
        n3895), .ZN(n571) );
  AOI222_X1 U426 ( .A1(Element[19]), .A2(n3927), .B1(\U52/DATA1_19 ), .B2(
        n3922), .C1(n3889), .C2(n573), .ZN(n572) );
  OAI222_X2 U427 ( .A1(n574), .A2(n3920), .B1(n3919), .B2(n4091), .C1(WireY), 
        .C2(n575), .ZN(n573) );
  OAI211_X2 U428 ( .C1(n3924), .C2(n4090), .A(n559), .B(n560), .ZN(n1052) );
  AOI22_X2 U429 ( .A1(\U95/DATA1_20 ), .A2(n3911), .B1(\U93/DATA1_20 ), .B2(
        n3895), .ZN(n559) );
  AOI222_X1 U430 ( .A1(Element[20]), .A2(n3927), .B1(\U52/DATA1_20 ), .B2(
        n3922), .C1(n3889), .C2(n561), .ZN(n560) );
  OAI222_X2 U432 ( .A1(n562), .A2(n3921), .B1(n3919), .B2(n4090), .C1(WireY), 
        .C2(n563), .ZN(n561) );
  OAI211_X2 U434 ( .C1(n3924), .C2(n4089), .A(n547), .B(n548), .ZN(n1051) );
  AOI22_X2 U436 ( .A1(\U95/DATA1_21 ), .A2(n3911), .B1(\U93/DATA1_21 ), .B2(
        n3895), .ZN(n547) );
  AOI222_X1 U437 ( .A1(Element[21]), .A2(n3927), .B1(\U52/DATA1_21 ), .B2(
        n3922), .C1(n3889), .C2(n549), .ZN(n548) );
  OAI222_X2 U438 ( .A1(n550), .A2(n3920), .B1(n3919), .B2(n4089), .C1(WireY), 
        .C2(n551), .ZN(n549) );
  OAI211_X2 U439 ( .C1(n3924), .C2(n4088), .A(n535), .B(n536), .ZN(n1050) );
  AOI22_X2 U440 ( .A1(\U95/DATA1_22 ), .A2(n3911), .B1(\U93/DATA1_22 ), .B2(
        n3895), .ZN(n535) );
  AOI222_X1 U441 ( .A1(Element[22]), .A2(n3927), .B1(\U52/DATA1_22 ), .B2(
        n3922), .C1(n3889), .C2(n537), .ZN(n536) );
  OAI222_X2 U442 ( .A1(n538), .A2(n3921), .B1(n3919), .B2(n4088), .C1(WireY), 
        .C2(n539), .ZN(n537) );
  OAI211_X2 U444 ( .C1(n3924), .C2(n4087), .A(n523), .B(n524), .ZN(n1049) );
  AOI22_X2 U446 ( .A1(\U95/DATA1_23 ), .A2(n3911), .B1(\U93/DATA1_23 ), .B2(
        n3895), .ZN(n523) );
  AOI222_X1 U448 ( .A1(Element[23]), .A2(n3927), .B1(\U52/DATA1_23 ), .B2(
        n3922), .C1(n3889), .C2(n525), .ZN(n524) );
  OAI222_X2 U449 ( .A1(n526), .A2(n3920), .B1(n3919), .B2(n4087), .C1(WireY), 
        .C2(n527), .ZN(n525) );
  OAI211_X2 U450 ( .C1(n3924), .C2(n4086), .A(n511), .B(n512), .ZN(n1048) );
  AOI22_X2 U451 ( .A1(\U95/DATA1_24 ), .A2(n3912), .B1(\U93/DATA1_24 ), .B2(
        n3895), .ZN(n511) );
  AOI222_X1 U452 ( .A1(Element[24]), .A2(n3927), .B1(\U52/DATA1_24 ), .B2(n215), .C1(n3889), .C2(n513), .ZN(n512) );
  OAI222_X2 U453 ( .A1(n514), .A2(n3920), .B1(n3919), .B2(n4086), .C1(WireY), 
        .C2(n515), .ZN(n513) );
  OAI211_X2 U454 ( .C1(n3924), .C2(n4085), .A(n499), .B(n500), .ZN(n1047) );
  AOI22_X2 U456 ( .A1(\U95/DATA1_25 ), .A2(n3912), .B1(\U93/DATA1_25 ), .B2(
        n3895), .ZN(n499) );
  AOI222_X1 U458 ( .A1(Element[25]), .A2(n3927), .B1(\U52/DATA1_25 ), .B2(n215), .C1(n3889), .C2(n501), .ZN(n500) );
  OAI222_X2 U460 ( .A1(n502), .A2(n3920), .B1(n3919), .B2(n4085), .C1(WireY), 
        .C2(n503), .ZN(n501) );
  OAI211_X2 U461 ( .C1(n3924), .C2(n4084), .A(n487), .B(n488), .ZN(n1046) );
  AOI22_X2 U462 ( .A1(\U95/DATA1_26 ), .A2(n3912), .B1(\U93/DATA1_26 ), .B2(
        n3895), .ZN(n487) );
  AOI222_X1 U463 ( .A1(Element[26]), .A2(n3927), .B1(\U52/DATA1_26 ), .B2(n215), .C1(n3889), .C2(n489), .ZN(n488) );
  OAI222_X2 U464 ( .A1(n490), .A2(n3920), .B1(n3919), .B2(n4084), .C1(WireY), 
        .C2(n491), .ZN(n489) );
  OAI211_X2 U465 ( .C1(n3924), .C2(n4083), .A(n475), .B(n476), .ZN(n1045) );
  AOI22_X2 U466 ( .A1(\U95/DATA1_27 ), .A2(n3912), .B1(\U93/DATA1_27 ), .B2(
        n3895), .ZN(n475) );
  AOI222_X1 U468 ( .A1(Element[27]), .A2(n3927), .B1(\U52/DATA1_27 ), .B2(n215), .C1(n3889), .C2(n477), .ZN(n476) );
  OAI222_X2 U470 ( .A1(n478), .A2(n3920), .B1(n3919), .B2(n4083), .C1(WireY), 
        .C2(n479), .ZN(n477) );
  OAI211_X2 U472 ( .C1(n3924), .C2(n4082), .A(n463), .B(n464), .ZN(n1044) );
  AOI22_X2 U473 ( .A1(\U95/DATA1_28 ), .A2(n3912), .B1(\U93/DATA1_28 ), .B2(
        n3895), .ZN(n463) );
  AOI222_X1 U474 ( .A1(Element[28]), .A2(n3927), .B1(\U52/DATA1_28 ), .B2(n215), .C1(n3889), .C2(n465), .ZN(n464) );
  OAI222_X2 U475 ( .A1(n466), .A2(n3920), .B1(n3919), .B2(n4082), .C1(WireY), 
        .C2(n467), .ZN(n465) );
  OAI211_X2 U476 ( .C1(n3924), .C2(n4081), .A(n451), .B(n452), .ZN(n1043) );
  AOI22_X2 U477 ( .A1(\U95/DATA1_29 ), .A2(n3912), .B1(\U93/DATA1_29 ), .B2(
        n3895), .ZN(n451) );
  AOI222_X1 U478 ( .A1(Element[29]), .A2(n3927), .B1(\U52/DATA1_29 ), .B2(n215), .C1(n3889), .C2(n453), .ZN(n452) );
  OAI222_X2 U480 ( .A1(n454), .A2(n3920), .B1(n3919), .B2(n4081), .C1(WireY), 
        .C2(n455), .ZN(n453) );
  OAI211_X2 U482 ( .C1(n3924), .C2(n4080), .A(n439), .B(n440), .ZN(n1042) );
  AOI22_X2 U484 ( .A1(\U95/DATA1_30 ), .A2(n3912), .B1(\U93/DATA1_30 ), .B2(
        n3895), .ZN(n439) );
  AOI222_X1 U485 ( .A1(Element[30]), .A2(n3927), .B1(\U52/DATA1_30 ), .B2(n215), .C1(n3889), .C2(n441), .ZN(n440) );
  OAI222_X2 U486 ( .A1(n442), .A2(n3920), .B1(n3919), .B2(n4080), .C1(WireY), 
        .C2(n443), .ZN(n441) );
  OAI211_X2 U487 ( .C1(n3924), .C2(n4079), .A(n427), .B(n428), .ZN(n1041) );
  AOI22_X2 U488 ( .A1(\U95/DATA1_31 ), .A2(n3912), .B1(\U93/DATA1_31 ), .B2(
        n3895), .ZN(n427) );
  AOI222_X1 U489 ( .A1(Element[31]), .A2(n3927), .B1(\U52/DATA1_31 ), .B2(n215), .C1(n3889), .C2(n429), .ZN(n428) );
  OAI222_X2 U490 ( .A1(n430), .A2(n3920), .B1(n3919), .B2(n4079), .C1(WireY), 
        .C2(n431), .ZN(n429) );
  OAI211_X2 U492 ( .C1(n212), .C2(n4078), .A(n415), .B(n416), .ZN(n1040) );
  AOI22_X2 U494 ( .A1(\U95/DATA1_32 ), .A2(n3912), .B1(\U93/DATA1_32 ), .B2(
        n3895), .ZN(n415) );
  AOI222_X1 U496 ( .A1(Element[32]), .A2(n3927), .B1(\U52/DATA1_32 ), .B2(n215), .C1(n3889), .C2(n417), .ZN(n416) );
  OAI222_X2 U497 ( .A1(n418), .A2(n3920), .B1(n3919), .B2(n4078), .C1(WireY), 
        .C2(n419), .ZN(n417) );
  OAI211_X2 U498 ( .C1(n212), .C2(n4077), .A(n403), .B(n404), .ZN(n1039) );
  AOI22_X2 U499 ( .A1(\U95/DATA1_33 ), .A2(n3912), .B1(\U93/DATA1_33 ), .B2(
        n3895), .ZN(n403) );
  AOI222_X1 U500 ( .A1(Element[33]), .A2(n3927), .B1(\U52/DATA1_33 ), .B2(n215), .C1(n3889), .C2(n405), .ZN(n404) );
  OAI222_X2 U501 ( .A1(n406), .A2(n3920), .B1(n3919), .B2(n4077), .C1(WireY), 
        .C2(n407), .ZN(n405) );
  OAI211_X2 U502 ( .C1(n212), .C2(n4076), .A(n391), .B(n392), .ZN(n1038) );
  AOI22_X2 U504 ( .A1(\U95/DATA1_34 ), .A2(n3912), .B1(\U93/DATA1_34 ), .B2(
        n3895), .ZN(n391) );
  AOI222_X1 U506 ( .A1(Element[34]), .A2(n3927), .B1(\U52/DATA1_34 ), .B2(n215), .C1(n3889), .C2(n393), .ZN(n392) );
  OAI222_X2 U508 ( .A1(n394), .A2(n3920), .B1(n3919), .B2(n4076), .C1(n3908), 
        .C2(n395), .ZN(n393) );
  OAI211_X2 U509 ( .C1(n3924), .C2(n4075), .A(n379), .B(n380), .ZN(n1037) );
  AOI22_X2 U510 ( .A1(\U95/DATA1_35 ), .A2(n3912), .B1(\U93/DATA1_35 ), .B2(
        n3895), .ZN(n379) );
  AOI222_X1 U511 ( .A1(Element[35]), .A2(n3927), .B1(\U52/DATA1_35 ), .B2(n215), .C1(n3889), .C2(n381), .ZN(n380) );
  OAI222_X2 U512 ( .A1(n382), .A2(n3920), .B1(n3919), .B2(n4075), .C1(n3908), 
        .C2(n383), .ZN(n381) );
  OAI211_X2 U513 ( .C1(n212), .C2(n4110), .A(n799), .B(n800), .ZN(n1072) );
  AOI22_X2 U514 ( .A1(\U95/DATA1_0 ), .A2(n3911), .B1(\U93/DATA1_0 ), .B2(
        n3895), .ZN(n799) );
  AOI222_X1 U516 ( .A1(Element[0]), .A2(n3927), .B1(\U52/DATA1_0 ), .B2(n3922), 
        .C1(n3889), .C2(n801), .ZN(n800) );
  OAI222_X2 U518 ( .A1(n802), .A2(n3921), .B1(n3919), .B2(n4110), .C1(WireY), 
        .C2(n803), .ZN(n801) );
  OAI211_X2 U520 ( .C1(n212), .C2(n4109), .A(n787), .B(n788), .ZN(n1071) );
  AOI22_X2 U521 ( .A1(\U95/DATA1_1 ), .A2(n3912), .B1(\U93/DATA1_1 ), .B2(
        n3895), .ZN(n787) );
  AOI222_X1 U522 ( .A1(Element[1]), .A2(n3927), .B1(\U52/DATA1_1 ), .B2(n215), 
        .C1(n3889), .C2(n789), .ZN(n788) );
  OAI222_X2 U523 ( .A1(n790), .A2(n3921), .B1(n3919), .B2(n4109), .C1(WireY), 
        .C2(n791), .ZN(n789) );
  OAI211_X2 U524 ( .C1(n212), .C2(n4108), .A(n775), .B(n776), .ZN(n1070) );
  AOI22_X2 U525 ( .A1(\U95/DATA1_2 ), .A2(n3912), .B1(\U93/DATA1_2 ), .B2(
        n3895), .ZN(n775) );
  AOI222_X1 U526 ( .A1(Element[2]), .A2(n3927), .B1(\U52/DATA1_2 ), .B2(n215), 
        .C1(n3889), .C2(n777), .ZN(n776) );
  OAI222_X2 U528 ( .A1(n778), .A2(n3921), .B1(n3919), .B2(n4108), .C1(WireY), 
        .C2(n779), .ZN(n777) );
  OAI211_X2 U530 ( .C1(n212), .C2(n4107), .A(n763), .B(n764), .ZN(n1069) );
  AOI22_X2 U532 ( .A1(\U95/DATA1_3 ), .A2(n3911), .B1(\U93/DATA1_3 ), .B2(
        n3895), .ZN(n763) );
  AOI222_X1 U533 ( .A1(Element[3]), .A2(n3927), .B1(\U52/DATA1_3 ), .B2(n215), 
        .C1(n3889), .C2(n765), .ZN(n764) );
  OAI222_X2 U534 ( .A1(n766), .A2(n3921), .B1(n3919), .B2(n4107), .C1(n3908), 
        .C2(n767), .ZN(n765) );
  OAI211_X2 U535 ( .C1(n212), .C2(n4106), .A(n751), .B(n752), .ZN(n1068) );
  AOI22_X2 U536 ( .A1(\U95/DATA1_4 ), .A2(n3912), .B1(\U93/DATA1_4 ), .B2(
        n3895), .ZN(n751) );
  AOI222_X1 U537 ( .A1(Element[4]), .A2(n3927), .B1(\U52/DATA1_4 ), .B2(n215), 
        .C1(n3889), .C2(n753), .ZN(n752) );
  OAI222_X2 U538 ( .A1(n754), .A2(n3921), .B1(n3919), .B2(n4106), .C1(WireY), 
        .C2(n755), .ZN(n753) );
  OAI211_X2 U540 ( .C1(n212), .C2(n4105), .A(n739), .B(n740), .ZN(n1067) );
  AOI22_X2 U542 ( .A1(\U95/DATA1_5 ), .A2(n3911), .B1(\U93/DATA1_5 ), .B2(
        n3895), .ZN(n739) );
  AOI222_X1 U544 ( .A1(Element[5]), .A2(n3927), .B1(\U52/DATA1_5 ), .B2(n215), 
        .C1(n3889), .C2(n741), .ZN(n740) );
  OAI222_X2 U545 ( .A1(n742), .A2(n3921), .B1(n3919), .B2(n4105), .C1(WireY), 
        .C2(n743), .ZN(n741) );
  OAI211_X2 U546 ( .C1(n212), .C2(n4104), .A(n727), .B(n728), .ZN(n1066) );
  AOI22_X2 U547 ( .A1(\U95/DATA1_6 ), .A2(n3911), .B1(\U93/DATA1_6 ), .B2(
        n3895), .ZN(n727) );
  AOI222_X1 U548 ( .A1(Element[6]), .A2(n3927), .B1(\U52/DATA1_6 ), .B2(n215), 
        .C1(n3889), .C2(n729), .ZN(n728) );
  OAI222_X2 U549 ( .A1(n730), .A2(n3921), .B1(n3919), .B2(n4104), .C1(n3908), 
        .C2(n731), .ZN(n729) );
  OAI211_X2 U550 ( .C1(n212), .C2(n4103), .A(n715), .B(n716), .ZN(n1065) );
  AOI22_X2 U552 ( .A1(\U95/DATA1_7 ), .A2(n3912), .B1(\U93/DATA1_7 ), .B2(
        n3895), .ZN(n715) );
  AOI222_X1 U554 ( .A1(Element[7]), .A2(n3927), .B1(\U52/DATA1_7 ), .B2(n215), 
        .C1(n3889), .C2(n717), .ZN(n716) );
  OAI222_X2 U556 ( .A1(n718), .A2(n3921), .B1(n3919), .B2(n4103), .C1(WireY), 
        .C2(n719), .ZN(n717) );
  OAI211_X2 U557 ( .C1(n212), .C2(n4102), .A(n703), .B(n704), .ZN(n1064) );
  AOI22_X2 U558 ( .A1(\U95/DATA1_8 ), .A2(n3912), .B1(\U93/DATA1_8 ), .B2(
        n3895), .ZN(n703) );
  AOI222_X1 U559 ( .A1(Element[8]), .A2(n3927), .B1(\U52/DATA1_8 ), .B2(n215), 
        .C1(n3889), .C2(n705), .ZN(n704) );
  OAI222_X2 U560 ( .A1(n706), .A2(n3921), .B1(n3919), .B2(n4102), .C1(WireY), 
        .C2(n707), .ZN(n705) );
  OAI211_X2 U561 ( .C1(n3924), .C2(n4101), .A(n691), .B(n692), .ZN(n1063) );
  AOI22_X2 U562 ( .A1(\U95/DATA1_9 ), .A2(n3911), .B1(\U93/DATA1_9 ), .B2(
        n3895), .ZN(n691) );
  AOI222_X1 U564 ( .A1(Element[9]), .A2(n3927), .B1(\U52/DATA1_9 ), .B2(n3922), 
        .C1(n3889), .C2(n693), .ZN(n692) );
  OAI222_X2 U566 ( .A1(n694), .A2(n3921), .B1(n3919), .B2(n4101), .C1(WireY), 
        .C2(n695), .ZN(n693) );
  OAI211_X2 U568 ( .C1(n3924), .C2(n4100), .A(n679), .B(n680), .ZN(n1062) );
  AOI22_X2 U569 ( .A1(\U95/DATA1_10 ), .A2(n3912), .B1(\U93/DATA1_10 ), .B2(
        n3895), .ZN(n679) );
  AOI222_X1 U570 ( .A1(Element[10]), .A2(n3927), .B1(\U52/DATA1_10 ), .B2(
        n3922), .C1(n3889), .C2(n681), .ZN(n680) );
  OAI222_X2 U571 ( .A1(n682), .A2(n3921), .B1(n3919), .B2(n4100), .C1(WireY), 
        .C2(n683), .ZN(n681) );
  OAI211_X2 U572 ( .C1(n3924), .C2(n4099), .A(n667), .B(n668), .ZN(n1061) );
  AOI22_X2 U573 ( .A1(\U95/DATA1_11 ), .A2(n3911), .B1(\U93/DATA1_11 ), .B2(
        n3895), .ZN(n667) );
  AOI222_X1 U574 ( .A1(Element[11]), .A2(n3927), .B1(\U52/DATA1_11 ), .B2(
        n3922), .C1(n3889), .C2(n669), .ZN(n668) );
  OAI222_X2 U576 ( .A1(n670), .A2(n3921), .B1(n3919), .B2(n4099), .C1(WireY), 
        .C2(n671), .ZN(n669) );
  OAI211_X2 U578 ( .C1(n3924), .C2(n4074), .A(n367), .B(n368), .ZN(n1036) );
  AOI22_X2 U580 ( .A1(\U95/DATA1_36 ), .A2(n3912), .B1(\U93/DATA1_36 ), .B2(
        n3895), .ZN(n367) );
  AOI222_X1 U581 ( .A1(Element[36]), .A2(n3927), .B1(\U52/DATA1_36 ), .B2(
        n3922), .C1(n3889), .C2(n369), .ZN(n368) );
  OAI222_X2 U582 ( .A1(n370), .A2(n3920), .B1(n3919), .B2(n4074), .C1(n3908), 
        .C2(n371), .ZN(n369) );
  OAI211_X2 U583 ( .C1(n3924), .C2(n4073), .A(n355), .B(n356), .ZN(n1035) );
  AOI22_X2 U584 ( .A1(\U95/DATA1_37 ), .A2(n3911), .B1(\U93/DATA1_37 ), .B2(
        n3895), .ZN(n355) );
  AOI222_X1 U585 ( .A1(Element[37]), .A2(n3927), .B1(\U52/DATA1_37 ), .B2(
        n3922), .C1(n3889), .C2(n357), .ZN(n356) );
  OAI222_X2 U586 ( .A1(n358), .A2(n3921), .B1(n3919), .B2(n4073), .C1(n3908), 
        .C2(n359), .ZN(n357) );
  OAI211_X2 U589 ( .C1(n3924), .C2(n4072), .A(n343), .B(n344), .ZN(n1034) );
  AOI22_X2 U591 ( .A1(\U95/DATA1_38 ), .A2(n3912), .B1(\U93/DATA1_38 ), .B2(
        n3895), .ZN(n343) );
  AOI222_X1 U592 ( .A1(Element[38]), .A2(n3927), .B1(\U52/DATA1_38 ), .B2(
        n3922), .C1(n3889), .C2(n345), .ZN(n344) );
  OAI222_X2 U594 ( .A1(n346), .A2(n3920), .B1(n3919), .B2(n4072), .C1(n3908), 
        .C2(n347), .ZN(n345) );
  OAI211_X2 U595 ( .C1(n3924), .C2(n4071), .A(n331), .B(n332), .ZN(n1033) );
  AOI22_X2 U596 ( .A1(\U95/DATA1_39 ), .A2(n3911), .B1(\U93/DATA1_39 ), .B2(
        n3895), .ZN(n331) );
  AOI222_X1 U598 ( .A1(Element[39]), .A2(n3927), .B1(\U52/DATA1_39 ), .B2(n215), .C1(n3889), .C2(n333), .ZN(n332) );
  OAI222_X2 U599 ( .A1(n334), .A2(n3921), .B1(n3919), .B2(n4071), .C1(n3908), 
        .C2(n335), .ZN(n333) );
  OAI211_X2 U604 ( .C1(n3924), .C2(n4070), .A(n319), .B(n320), .ZN(n1032) );
  AOI22_X2 U606 ( .A1(\U95/DATA1_40 ), .A2(n3912), .B1(\U93/DATA1_40 ), .B2(
        n3895), .ZN(n319) );
  AOI222_X1 U607 ( .A1(Element[40]), .A2(n3927), .B1(\U52/DATA1_40 ), .B2(n215), .C1(n3889), .C2(n321), .ZN(n320) );
  OAI222_X2 U609 ( .A1(n322), .A2(n3921), .B1(n3919), .B2(n4070), .C1(n3908), 
        .C2(n323), .ZN(n321) );
  OAI211_X2 U610 ( .C1(n3924), .C2(n4069), .A(n307), .B(n308), .ZN(n1031) );
  AOI22_X2 U614 ( .A1(\U95/DATA1_41 ), .A2(n3911), .B1(\U93/DATA1_41 ), .B2(
        n3895), .ZN(n307) );
  AOI222_X1 U618 ( .A1(Element[41]), .A2(n3927), .B1(\U52/DATA1_41 ), .B2(n215), .C1(n3889), .C2(n309), .ZN(n308) );
  OAI222_X2 U706 ( .A1(n310), .A2(n3920), .B1(n3919), .B2(n4069), .C1(n3908), 
        .C2(n311), .ZN(n309) );
  OAI211_X2 U708 ( .C1(n3924), .C2(n4068), .A(n295), .B(n296), .ZN(n1030) );
  AOI22_X2 U709 ( .A1(\U95/DATA1_42 ), .A2(n3912), .B1(\U93/DATA1_42 ), .B2(
        n3895), .ZN(n295) );
  AOI222_X1 U713 ( .A1(Element[42]), .A2(n3927), .B1(\U52/DATA1_42 ), .B2(n215), .C1(n3889), .C2(n297), .ZN(n296) );
  OAI222_X2 U714 ( .A1(n298), .A2(n3920), .B1(n220), .B2(n4068), .C1(n3908), 
        .C2(n299), .ZN(n297) );
  OAI211_X2 U715 ( .C1(n3924), .C2(n4067), .A(n283), .B(n284), .ZN(n1029) );
  AOI22_X2 U716 ( .A1(\U95/DATA1_43 ), .A2(n3911), .B1(\U93/DATA1_43 ), .B2(
        n3895), .ZN(n283) );
  AOI222_X1 U717 ( .A1(Element[43]), .A2(n3927), .B1(\U52/DATA1_43 ), .B2(n215), .C1(n3889), .C2(n285), .ZN(n284) );
  OAI222_X2 U718 ( .A1(n286), .A2(n3921), .B1(n3919), .B2(n4067), .C1(n3908), 
        .C2(n287), .ZN(n285) );
  OAI211_X2 U719 ( .C1(n3924), .C2(n4066), .A(n271), .B(n272), .ZN(n1028) );
  AOI22_X2 U720 ( .A1(\U95/DATA1_44 ), .A2(n3912), .B1(\U93/DATA1_44 ), .B2(
        n3895), .ZN(n271) );
  AOI222_X1 U721 ( .A1(Element[44]), .A2(n3927), .B1(\U52/DATA1_44 ), .B2(n215), .C1(n3889), .C2(n273), .ZN(n272) );
  OAI222_X2 U722 ( .A1(n274), .A2(n3920), .B1(n220), .B2(n4066), .C1(n3908), 
        .C2(n275), .ZN(n273) );
  OAI211_X2 U723 ( .C1(n3924), .C2(n4065), .A(n259), .B(n260), .ZN(n1027) );
  AOI22_X2 U724 ( .A1(\U95/DATA1_45 ), .A2(n3911), .B1(\U93/DATA1_45 ), .B2(
        n3895), .ZN(n259) );
  AOI222_X1 U725 ( .A1(Element[45]), .A2(n3927), .B1(\U52/DATA1_45 ), .B2(n215), .C1(n3889), .C2(n261), .ZN(n260) );
  OAI222_X2 U728 ( .A1(n262), .A2(n3921), .B1(n3919), .B2(n4065), .C1(n3908), 
        .C2(n263), .ZN(n261) );
  OAI211_X2 U730 ( .C1(n3924), .C2(n4064), .A(n247), .B(n248), .ZN(n1026) );
  AOI22_X2 U734 ( .A1(\U95/DATA1_46 ), .A2(n3912), .B1(\U93/DATA1_46 ), .B2(
        n3895), .ZN(n247) );
  AOI222_X1 U823 ( .A1(Element[46]), .A2(n3927), .B1(\U52/DATA1_46 ), .B2(n215), .C1(n3889), .C2(n249), .ZN(n248) );
  OAI222_X2 U825 ( .A1(n250), .A2(n3921), .B1(n220), .B2(n4064), .C1(n3908), 
        .C2(n251), .ZN(n249) );
  OAI211_X2 U827 ( .C1(n3924), .C2(n4063), .A(n213), .B(n214), .ZN(n1025) );
  AOI22_X2 U828 ( .A1(\U95/DATA1_47 ), .A2(n3911), .B1(\U93/DATA1_47 ), .B2(
        n3895), .ZN(n213) );
  AOI222_X1 U829 ( .A1(Element[47]), .A2(n3927), .B1(\U52/DATA1_47 ), .B2(n215), .C1(n3889), .C2(n217), .ZN(n214) );
  OAI222_X2 U830 ( .A1(n218), .A2(n3920), .B1(n4063), .B2(n3919), .C1(WireY), 
        .C2(n221), .ZN(n217) );
  AOI22_X2 U831 ( .A1(PosRowY[11]), .A2(n921), .B1(Row_noY[9]), .B2(n3907), 
        .ZN(n936) );
  AOI22_X2 U832 ( .A1(PosRowY[10]), .A2(n921), .B1(Row_noY[8]), .B2(n3907), 
        .ZN(n935) );
  AOI22_X2 U833 ( .A1(PosRowY[9]), .A2(n921), .B1(Row_noY[7]), .B2(n3907), 
        .ZN(n934) );
  AOI22_X2 U834 ( .A1(PosRowY[8]), .A2(n921), .B1(Row_noY[6]), .B2(n3907), 
        .ZN(n933) );
  AOI22_X2 U835 ( .A1(PosRowY[7]), .A2(n921), .B1(Row_noY[5]), .B2(n3907), 
        .ZN(n932) );
  AOI22_X2 U836 ( .A1(PosRowY[6]), .A2(n921), .B1(Row_noY[4]), .B2(n3907), 
        .ZN(n931) );
  AOI22_X2 U837 ( .A1(PosRowY[5]), .A2(n921), .B1(Row_noY[3]), .B2(n3907), 
        .ZN(n930) );
  AOI22_X2 U838 ( .A1(PosRowY[4]), .A2(n921), .B1(Row_noY[2]), .B2(n3907), 
        .ZN(n929) );
  AOI22_X2 U839 ( .A1(PosRowY[3]), .A2(n921), .B1(Row_noY[1]), .B2(n3907), 
        .ZN(n928) );
  OAI21_X2 U840 ( .B1(n835), .B2(n35), .A(n3953), .ZN(n1073) );
  OAI21_X2 U841 ( .B1(n938), .B2(n28), .A(n921), .ZN(n1077) );
  OAI21_X2 U842 ( .B1(n920), .B2(n921), .A(n922), .ZN(n1075) );
  OAI21_X2 U843 ( .B1(n193), .B2(n3953), .A(n194), .ZN(n1023) );
  AOI22_X2 U844 ( .A1(PosRowX[11]), .A2(n3953), .B1(Row_noX[9]), .B2(n201), 
        .ZN(n210) );
  AOI22_X2 U845 ( .A1(PosRowX[10]), .A2(n3953), .B1(Row_noX[8]), .B2(n201), 
        .ZN(n209) );
  AOI22_X2 U846 ( .A1(PosRowX[9]), .A2(n3953), .B1(Row_noX[7]), .B2(n201), 
        .ZN(n208) );
  AOI22_X2 U847 ( .A1(PosRowX[8]), .A2(n3953), .B1(Row_noX[6]), .B2(n201), 
        .ZN(n207) );
  AOI22_X2 U848 ( .A1(PosRowX[7]), .A2(n3953), .B1(Row_noX[5]), .B2(n201), 
        .ZN(n206) );
  AOI22_X2 U849 ( .A1(PosRowX[6]), .A2(n3953), .B1(Row_noX[4]), .B2(n201), 
        .ZN(n205) );
  AOI22_X2 U850 ( .A1(PosRowX[5]), .A2(n3953), .B1(Row_noX[3]), .B2(n201), 
        .ZN(n204) );
  AOI22_X2 U851 ( .A1(PosRowX[4]), .A2(n3953), .B1(Row_noX[2]), .B2(n201), 
        .ZN(n203) );
  AOI22_X2 U852 ( .A1(PosRowX[3]), .A2(n3953), .B1(Row_noX[1]), .B2(n201), 
        .ZN(n202) );
  AOI22_X2 U853 ( .A1(PosRowX[2]), .A2(n3953), .B1(Row_noX[0]), .B2(n201), 
        .ZN(n200) );
  AOI22_X2 U854 ( .A1(PosRowY[2]), .A2(n921), .B1(Row_noY[0]), .B2(n3907), 
        .ZN(n927) );
  AOI22_X2 U855 ( .A1(PosRowY[12]), .A2(n921), .B1(Row_noY[10]), .B2(n3907), 
        .ZN(n937) );
  AOI22_X2 U856 ( .A1(PosRowX[12]), .A2(n3953), .B1(Row_noX[10]), .B2(n201), 
        .ZN(n211) );
  INV_X4 U857 ( .A(n824), .ZN(n3927) );
  INV_X4 U858 ( .A(n927), .ZN(n3928) );
  INV_X4 U859 ( .A(n928), .ZN(n3929) );
  INV_X4 U860 ( .A(n929), .ZN(n3930) );
  INV_X4 U861 ( .A(n930), .ZN(n3931) );
  INV_X4 U862 ( .A(n931), .ZN(n3932) );
  INV_X4 U863 ( .A(n932), .ZN(n3933) );
  INV_X4 U864 ( .A(n933), .ZN(n3934) );
  INV_X4 U865 ( .A(n934), .ZN(n3935) );
  INV_X4 U866 ( .A(n935), .ZN(n3936) );
  INV_X4 U867 ( .A(n936), .ZN(n3937) );
  INV_X4 U868 ( .A(n937), .ZN(n3938) );
  INV_X4 U869 ( .A(n827), .ZN(n3939) );
  INV_X4 U870 ( .A(n818), .ZN(n3940) );
  INV_X4 U871 ( .A(n836), .ZN(WireX) );
  INV_X4 U872 ( .A(n200), .ZN(n3942) );
  INV_X4 U873 ( .A(n202), .ZN(n3943) );
  INV_X4 U874 ( .A(n203), .ZN(n3944) );
  INV_X4 U875 ( .A(n204), .ZN(n3945) );
  INV_X4 U876 ( .A(n205), .ZN(n3946) );
  INV_X4 U877 ( .A(n206), .ZN(n3947) );
  INV_X4 U878 ( .A(n207), .ZN(n3948) );
  INV_X4 U879 ( .A(n208), .ZN(n3949) );
  INV_X4 U880 ( .A(n209), .ZN(n3950) );
  INV_X4 U881 ( .A(n210), .ZN(n3951) );
  INV_X4 U882 ( .A(n211), .ZN(n3952) );
  INV_X4 U883 ( .A(n819), .ZN(n3954) );
  INV_X4 U884 ( .A(n837), .ZN(n3955) );
  INV_X4 U885 ( .A(PosDX[0]), .ZN(n3956) );
  INV_X4 U886 ( .A(n941), .ZN(n3957) );
  INV_X4 U887 ( .A(PosDY[0]), .ZN(n3958) );
  INV_X4 U888 ( .A(n832), .ZN(n3959) );
  INV_X4 U889 ( .A(n826), .ZN(n3960) );
  INV_X4 U890 ( .A(n920), .ZN(n3961) );
  INV_X4 U891 ( .A(n833), .ZN(n3962) );
  INV_X4 U892 ( .A(n926), .ZN(n3963) );
  INV_X4 U893 ( .A(n821), .ZN(n3964) );
  INV_X4 U894 ( .A(n193), .ZN(n3965) );
  INV_X4 U895 ( .A(n822), .ZN(n3966) );
  INV_X4 U896 ( .A(\U166/DATA1_47 ), .ZN(n3967) );
  INV_X4 U897 ( .A(\U166/DATA1_46 ), .ZN(n3968) );
  INV_X4 U898 ( .A(\U166/DATA1_45 ), .ZN(n3969) );
  INV_X4 U899 ( .A(\U166/DATA1_44 ), .ZN(n3970) );
  INV_X4 U900 ( .A(\U166/DATA1_43 ), .ZN(n3971) );
  INV_X4 U901 ( .A(\U166/DATA1_42 ), .ZN(n3972) );
  INV_X4 U902 ( .A(\U166/DATA1_41 ), .ZN(n3973) );
  INV_X4 U903 ( .A(\U166/DATA1_40 ), .ZN(n3974) );
  INV_X4 U904 ( .A(\U166/DATA1_39 ), .ZN(n3975) );
  INV_X4 U905 ( .A(\U166/DATA1_38 ), .ZN(n3976) );
  INV_X4 U906 ( .A(\U166/DATA1_37 ), .ZN(n3977) );
  INV_X4 U907 ( .A(\U166/DATA1_36 ), .ZN(n3978) );
  INV_X4 U908 ( .A(\U166/DATA1_35 ), .ZN(n3979) );
  INV_X4 U909 ( .A(\U166/DATA1_34 ), .ZN(n3980) );
  INV_X4 U910 ( .A(\U166/DATA1_33 ), .ZN(n3981) );
  INV_X4 U911 ( .A(\U166/DATA1_32 ), .ZN(n3982) );
  INV_X4 U912 ( .A(\U166/DATA1_31 ), .ZN(n3983) );
  INV_X4 U913 ( .A(\U166/DATA1_30 ), .ZN(n3984) );
  INV_X4 U914 ( .A(\U166/DATA1_29 ), .ZN(n3985) );
  INV_X4 U915 ( .A(\U166/DATA1_28 ), .ZN(n3986) );
  INV_X4 U916 ( .A(\U166/DATA1_27 ), .ZN(n3987) );
  INV_X4 U917 ( .A(\U166/DATA1_26 ), .ZN(n3988) );
  INV_X4 U918 ( .A(\U166/DATA1_25 ), .ZN(n3989) );
  INV_X4 U919 ( .A(\U166/DATA1_24 ), .ZN(n3990) );
  INV_X4 U920 ( .A(\U166/DATA1_23 ), .ZN(n3991) );
  INV_X4 U921 ( .A(\U166/DATA1_22 ), .ZN(n3992) );
  INV_X4 U922 ( .A(\U166/DATA1_21 ), .ZN(n3993) );
  INV_X4 U923 ( .A(\U166/DATA1_20 ), .ZN(n3994) );
  INV_X4 U924 ( .A(\U166/DATA1_19 ), .ZN(n3995) );
  INV_X4 U925 ( .A(\U166/DATA1_18 ), .ZN(n3996) );
  INV_X4 U926 ( .A(\U166/DATA1_17 ), .ZN(n3997) );
  INV_X4 U927 ( .A(\U166/DATA1_16 ), .ZN(n3998) );
  INV_X4 U928 ( .A(\U166/DATA1_15 ), .ZN(n3999) );
  INV_X4 U929 ( .A(\U166/DATA1_14 ), .ZN(n4000) );
  INV_X4 U930 ( .A(\U166/DATA1_13 ), .ZN(n4001) );
  INV_X4 U931 ( .A(\U166/DATA1_12 ), .ZN(n4002) );
  INV_X4 U932 ( .A(\U166/DATA1_11 ), .ZN(n4003) );
  INV_X4 U933 ( .A(\U166/DATA1_10 ), .ZN(n4004) );
  INV_X4 U934 ( .A(\U166/DATA1_9 ), .ZN(n4005) );
  INV_X4 U935 ( .A(\U166/DATA1_8 ), .ZN(n4006) );
  INV_X4 U936 ( .A(\U166/DATA1_7 ), .ZN(n4007) );
  INV_X4 U937 ( .A(\U166/DATA1_6 ), .ZN(n4008) );
  INV_X4 U938 ( .A(\U166/DATA1_5 ), .ZN(n4009) );
  INV_X4 U939 ( .A(\U166/DATA1_4 ), .ZN(n4010) );
  INV_X4 U940 ( .A(\U166/DATA1_3 ), .ZN(n4011) );
  INV_X4 U941 ( .A(\U166/DATA1_2 ), .ZN(n4012) );
  INV_X4 U942 ( .A(\U166/DATA1_1 ), .ZN(n4013) );
  INV_X4 U943 ( .A(\U166/DATA1_0 ), .ZN(n4014) );
  INV_X4 U944 ( .A(\U163/DATA1_47 ), .ZN(n4015) );
  INV_X4 U945 ( .A(\U163/DATA1_46 ), .ZN(n4016) );
  INV_X4 U946 ( .A(\U163/DATA1_45 ), .ZN(n4017) );
  INV_X4 U947 ( .A(\U163/DATA1_44 ), .ZN(n4018) );
  INV_X4 U948 ( .A(\U163/DATA1_43 ), .ZN(n4019) );
  INV_X4 U949 ( .A(\U163/DATA1_42 ), .ZN(n4020) );
  INV_X4 U950 ( .A(\U163/DATA1_41 ), .ZN(n4021) );
  INV_X4 U951 ( .A(\U163/DATA1_40 ), .ZN(n4022) );
  INV_X4 U952 ( .A(\U163/DATA1_39 ), .ZN(n4023) );
  INV_X4 U953 ( .A(\U163/DATA1_38 ), .ZN(n4024) );
  INV_X4 U954 ( .A(\U163/DATA1_37 ), .ZN(n4025) );
  INV_X4 U955 ( .A(\U163/DATA1_36 ), .ZN(n4026) );
  INV_X4 U956 ( .A(\U163/DATA1_35 ), .ZN(n4027) );
  INV_X4 U957 ( .A(\U163/DATA1_34 ), .ZN(n4028) );
  INV_X4 U958 ( .A(\U163/DATA1_33 ), .ZN(n4029) );
  INV_X4 U959 ( .A(\U163/DATA1_32 ), .ZN(n4030) );
  INV_X4 U960 ( .A(\U163/DATA1_31 ), .ZN(n4031) );
  INV_X4 U961 ( .A(\U163/DATA1_30 ), .ZN(n4032) );
  INV_X4 U962 ( .A(\U163/DATA1_29 ), .ZN(n4033) );
  INV_X4 U963 ( .A(\U163/DATA1_28 ), .ZN(n4034) );
  INV_X4 U964 ( .A(\U163/DATA1_27 ), .ZN(n4035) );
  INV_X4 U965 ( .A(\U163/DATA1_26 ), .ZN(n4036) );
  INV_X4 U966 ( .A(\U163/DATA1_25 ), .ZN(n4037) );
  INV_X4 U967 ( .A(\U163/DATA1_24 ), .ZN(n4038) );
  INV_X4 U968 ( .A(\U163/DATA1_23 ), .ZN(n4039) );
  INV_X4 U969 ( .A(\U163/DATA1_22 ), .ZN(n4040) );
  INV_X4 U970 ( .A(\U163/DATA1_21 ), .ZN(n4041) );
  INV_X4 U971 ( .A(\U163/DATA1_20 ), .ZN(n4042) );
  INV_X4 U972 ( .A(\U163/DATA1_19 ), .ZN(n4043) );
  INV_X4 U973 ( .A(\U163/DATA1_18 ), .ZN(n4044) );
  INV_X4 U974 ( .A(\U163/DATA1_17 ), .ZN(n4045) );
  INV_X4 U975 ( .A(\U163/DATA1_16 ), .ZN(n4046) );
  INV_X4 U976 ( .A(\U163/DATA1_15 ), .ZN(n4047) );
  INV_X4 U977 ( .A(\U163/DATA1_14 ), .ZN(n4048) );
  INV_X4 U978 ( .A(\U163/DATA1_13 ), .ZN(n4049) );
  INV_X4 U979 ( .A(\U163/DATA1_12 ), .ZN(n4050) );
  INV_X4 U980 ( .A(\U163/DATA1_11 ), .ZN(n4051) );
  INV_X4 U981 ( .A(\U163/DATA1_10 ), .ZN(n4052) );
  INV_X4 U982 ( .A(\U163/DATA1_9 ), .ZN(n4053) );
  INV_X4 U983 ( .A(\U163/DATA1_8 ), .ZN(n4054) );
  INV_X4 U984 ( .A(\U163/DATA1_7 ), .ZN(n4055) );
  INV_X4 U985 ( .A(\U163/DATA1_6 ), .ZN(n4056) );
  INV_X4 U986 ( .A(\U163/DATA1_5 ), .ZN(n4057) );
  INV_X4 U987 ( .A(\U163/DATA1_4 ), .ZN(n4058) );
  INV_X4 U988 ( .A(\U163/DATA1_3 ), .ZN(n4059) );
  INV_X4 U989 ( .A(\U163/DATA1_2 ), .ZN(n4060) );
  INV_X4 U990 ( .A(\U163/DATA1_1 ), .ZN(n4061) );
  INV_X4 U991 ( .A(\U163/DATA1_0 ), .ZN(n4062) );
  INV_X4 U992 ( .A(\U90/DATA1_47 ), .ZN(n4063) );
  INV_X4 U993 ( .A(\U90/DATA1_46 ), .ZN(n4064) );
  INV_X4 U994 ( .A(\U90/DATA1_45 ), .ZN(n4065) );
  INV_X4 U995 ( .A(\U90/DATA1_44 ), .ZN(n4066) );
  INV_X4 U996 ( .A(\U90/DATA1_43 ), .ZN(n4067) );
  INV_X4 U997 ( .A(\U90/DATA1_42 ), .ZN(n4068) );
  INV_X4 U998 ( .A(\U90/DATA1_41 ), .ZN(n4069) );
  INV_X4 U999 ( .A(\U90/DATA1_40 ), .ZN(n4070) );
  INV_X4 U1000 ( .A(\U90/DATA1_39 ), .ZN(n4071) );
  INV_X4 U1001 ( .A(\U90/DATA1_38 ), .ZN(n4072) );
  INV_X4 U1002 ( .A(\U90/DATA1_37 ), .ZN(n4073) );
  INV_X4 U1003 ( .A(\U90/DATA1_36 ), .ZN(n4074) );
  INV_X4 U1004 ( .A(\U90/DATA1_35 ), .ZN(n4075) );
  INV_X4 U1005 ( .A(\U90/DATA1_34 ), .ZN(n4076) );
  INV_X4 U1006 ( .A(\U90/DATA1_33 ), .ZN(n4077) );
  INV_X4 U1007 ( .A(\U90/DATA1_32 ), .ZN(n4078) );
  INV_X4 U1008 ( .A(\U90/DATA1_31 ), .ZN(n4079) );
  INV_X4 U1009 ( .A(\U90/DATA1_30 ), .ZN(n4080) );
  INV_X4 U1010 ( .A(\U90/DATA1_29 ), .ZN(n4081) );
  INV_X4 U1011 ( .A(\U90/DATA1_28 ), .ZN(n4082) );
  INV_X4 U1012 ( .A(\U90/DATA1_27 ), .ZN(n4083) );
  INV_X4 U1013 ( .A(\U90/DATA1_26 ), .ZN(n4084) );
  INV_X4 U1014 ( .A(\U90/DATA1_25 ), .ZN(n4085) );
  INV_X4 U1062 ( .A(\U90/DATA1_24 ), .ZN(n4086) );
  INV_X4 U1063 ( .A(\U90/DATA1_23 ), .ZN(n4087) );
  INV_X4 U1064 ( .A(\U90/DATA1_22 ), .ZN(n4088) );
  INV_X4 U1065 ( .A(\U90/DATA1_21 ), .ZN(n4089) );
  INV_X4 U1067 ( .A(\U90/DATA1_20 ), .ZN(n4090) );
  INV_X4 U1068 ( .A(\U90/DATA1_19 ), .ZN(n4091) );
  INV_X4 U1069 ( .A(\U90/DATA1_18 ), .ZN(n4092) );
  INV_X4 U1070 ( .A(\U90/DATA1_17 ), .ZN(n4093) );
  INV_X4 U1071 ( .A(\U90/DATA1_16 ), .ZN(n4094) );
  INV_X4 U1072 ( .A(\U90/DATA1_15 ), .ZN(n4095) );
  INV_X4 U1073 ( .A(\U90/DATA1_14 ), .ZN(n4096) );
  INV_X4 U1074 ( .A(\U90/DATA1_13 ), .ZN(n4097) );
  INV_X4 U1075 ( .A(\U90/DATA1_12 ), .ZN(n4098) );
  INV_X4 U1079 ( .A(\U90/DATA1_11 ), .ZN(n4099) );
  INV_X4 U1080 ( .A(\U90/DATA1_10 ), .ZN(n4100) );
  INV_X4 U1081 ( .A(\U90/DATA1_9 ), .ZN(n4101) );
  INV_X4 U1082 ( .A(\U90/DATA1_8 ), .ZN(n4102) );
  INV_X4 U1083 ( .A(\U90/DATA1_7 ), .ZN(n4103) );
  INV_X4 U1084 ( .A(\U90/DATA1_6 ), .ZN(n4104) );
  INV_X4 U1085 ( .A(\U90/DATA1_5 ), .ZN(n4105) );
  INV_X4 U1086 ( .A(\U90/DATA1_4 ), .ZN(n4106) );
  INV_X4 U1087 ( .A(\U90/DATA1_3 ), .ZN(n4107) );
  INV_X4 U1088 ( .A(\U90/DATA1_2 ), .ZN(n4108) );
  INV_X4 U1089 ( .A(\U90/DATA1_1 ), .ZN(n4109) );
  INV_X4 U1090 ( .A(\U90/DATA1_0 ), .ZN(n4110) );
endmodule


module arithController ( clock, reset, DiagonalX, DiagonalY, Element, 
        NewElement, EnableChange, SubInput1, SubInput2, AddInput1, AddInput2, 
        NewDiagonalX, NewDiagonalY, SubOutput, AddOutput, DiagonalXDone, 
        DiagonalYDone );
  input [47:0] DiagonalX;
  input [47:0] DiagonalY;
  input [47:0] Element;
  input [47:0] NewElement;
  output [23:0] SubInput1;
  output [23:0] SubInput2;
  output [23:0] AddInput1;
  output [23:0] AddInput2;
  output [47:0] NewDiagonalX;
  output [47:0] NewDiagonalY;
  input [23:0] SubOutput;
  input [23:0] AddOutput;
  input clock, reset, EnableChange;
  output DiagonalXDone, DiagonalYDone;
  wire   \U3/U1/DATA2_1 , \U3/U1/DATA2_2 , \U3/U1/DATA2_3 , \U12/DATA2_0 ,
         \U12/DATA2_1 , \U12/DATA2_2 , \U12/DATA2_3 , \U12/DATA2_4 ,
         \U12/DATA2_5 , \U12/DATA2_6 , \U12/DATA2_7 , \U12/DATA2_8 ,
         \U12/DATA2_9 , \U12/DATA2_10 , \U12/DATA2_11 , \U12/DATA2_12 ,
         \U12/DATA2_13 , \U12/DATA2_14 , \U12/DATA2_15 , \U12/DATA2_16 ,
         \U12/DATA2_17 , \U12/DATA2_18 , \U12/DATA2_19 , \U12/DATA2_20 ,
         \U12/DATA2_21 , \U12/DATA2_22 , \U12/DATA2_23 , \U12/DATA1_0 ,
         \U12/DATA1_1 , \U12/DATA1_2 , \U12/DATA1_3 , \U12/DATA1_4 ,
         \U12/DATA1_5 , \U12/DATA1_6 , \U12/DATA1_7 , \U12/DATA1_8 ,
         \U12/DATA1_9 , \U12/DATA1_10 , \U12/DATA1_11 , \U12/DATA1_12 ,
         \U12/DATA1_13 , \U12/DATA1_14 , \U12/DATA1_15 , \U12/DATA1_16 ,
         \U12/DATA1_17 , \U12/DATA1_18 , \U12/DATA1_19 , \U12/DATA1_20 ,
         \U12/DATA1_21 , \U12/DATA1_22 , \U12/DATA1_23 , \U11/DATA2_0 ,
         \U11/DATA2_1 , \U11/DATA2_2 , \U11/DATA2_3 , \U11/DATA2_4 ,
         \U11/DATA2_5 , \U11/DATA2_6 , \U11/DATA2_7 , \U11/DATA2_8 ,
         \U11/DATA2_9 , \U11/DATA2_10 , \U11/DATA2_11 , \U11/DATA2_12 ,
         \U11/DATA2_13 , \U11/DATA2_14 , \U11/DATA2_15 , \U11/DATA2_16 ,
         \U11/DATA2_17 , \U11/DATA2_18 , \U11/DATA2_19 , \U11/DATA2_20 ,
         \U11/DATA2_21 , \U11/DATA2_22 , \U11/DATA2_23 , \U11/DATA1_0 ,
         \U11/DATA1_1 , \U11/DATA1_2 , \U11/DATA1_3 , \U11/DATA1_4 ,
         \U11/DATA1_5 , \U11/DATA1_6 , \U11/DATA1_7 , \U11/DATA1_8 ,
         \U11/DATA1_9 , \U11/DATA1_10 , \U11/DATA1_11 , \U11/DATA1_12 ,
         \U11/DATA1_13 , \U11/DATA1_14 , \U11/DATA1_15 , \U11/DATA1_16 ,
         \U11/DATA1_17 , \U11/DATA1_18 , \U11/DATA1_19 , \U11/DATA1_20 ,
         \U11/DATA1_21 , \U11/DATA1_22 , \U11/DATA1_23 , \U8/Z_0 , \U8/Z_1 ,
         \U8/Z_2 , \U8/Z_3 , \U8/Z_4 , \U8/Z_5 , \U8/Z_6 , \U8/Z_7 , \U8/Z_8 ,
         \U8/Z_9 , \U8/Z_10 , \U8/Z_11 , \U8/Z_12 , \U8/Z_13 , \U8/Z_14 ,
         \U8/Z_15 , \U8/Z_16 , \U8/Z_17 , \U8/Z_18 , \U8/Z_19 , \U8/Z_20 ,
         \U8/Z_21 , \U8/Z_22 , \U8/Z_23 , \U7/Z_0 , \U7/Z_1 , \U7/Z_2 ,
         \U7/Z_3 , \U7/Z_4 , \U7/Z_5 , \U7/Z_6 , \U7/Z_7 , \U7/Z_8 , \U7/Z_9 ,
         \U7/Z_10 , \U7/Z_11 , \U7/Z_12 , \U7/Z_13 , \U7/Z_14 , \U7/Z_15 ,
         \U7/Z_16 , \U7/Z_17 , \U7/Z_18 , \U7/Z_19 , \U7/Z_20 , \U7/Z_21 ,
         \U7/Z_22 , \U7/Z_23 , \U6/DATA2_0 , \U6/DATA2_1 , \U6/DATA2_2 ,
         \U6/DATA2_3 , \U6/DATA2_4 , \U6/DATA2_5 , \U6/DATA2_6 , \U6/DATA2_7 ,
         \U6/DATA2_8 , \U6/DATA2_9 , \U6/DATA2_10 , \U6/DATA2_11 ,
         \U6/DATA2_12 , \U6/DATA2_13 , \U6/DATA2_14 , \U6/DATA2_15 ,
         \U6/DATA2_16 , \U6/DATA2_17 , \U6/DATA2_18 , \U6/DATA2_19 ,
         \U6/DATA2_20 , \U6/DATA2_21 , \U6/DATA2_22 , \U6/DATA2_23 ,
         \U6/DATA1_0 , \U6/DATA1_1 , \U6/DATA1_2 , \U6/DATA1_3 , \U6/DATA1_4 ,
         \U6/DATA1_5 , \U6/DATA1_6 , \U6/DATA1_7 , \U6/DATA1_8 , \U6/DATA1_9 ,
         \U6/DATA1_10 , \U6/DATA1_11 , \U6/DATA1_12 , \U6/DATA1_13 ,
         \U6/DATA1_14 , \U6/DATA1_15 , \U6/DATA1_16 , \U6/DATA1_17 ,
         \U6/DATA1_18 , \U6/DATA1_19 , \U6/DATA1_20 , \U6/DATA1_21 ,
         \U6/DATA1_22 , \U6/DATA1_23 , \U5/DATA1_0 , \U5/DATA1_1 ,
         \U5/DATA1_2 , \U5/DATA1_3 , \U5/DATA1_4 , \U5/DATA1_5 , \U5/DATA1_6 ,
         \U5/DATA1_7 , \U5/DATA1_8 , \U5/DATA1_9 , \U5/DATA1_10 ,
         \U5/DATA1_11 , \U5/DATA1_12 , \U5/DATA1_13 , \U5/DATA1_14 ,
         \U5/DATA1_15 , \U5/DATA1_16 , \U5/DATA1_17 , \U5/DATA1_18 ,
         \U5/DATA1_19 , \U5/DATA1_20 , \U5/DATA1_21 , \U5/DATA1_22 ,
         \U5/DATA1_23 , \U4/Z_0 , \U4/Z_1 , \U4/Z_2 , \U4/Z_3 , \U4/Z_4 ,
         \U4/Z_5 , \U4/Z_6 , \U4/Z_7 , \U4/Z_8 , \U4/Z_9 , \U4/Z_10 ,
         \U4/Z_11 , \U4/Z_12 , \U4/Z_13 , \U4/Z_14 , \U4/Z_15 , \U4/Z_16 ,
         \U4/Z_17 , \U4/Z_18 , \U4/Z_19 , \U4/Z_20 , \U4/Z_21 , \U4/Z_22 ,
         \U4/Z_23 , \U4/DATA1_0 , \U4/DATA1_1 , \U4/DATA1_2 , \U4/DATA1_3 ,
         \U4/DATA1_4 , \U4/DATA1_5 , \U4/DATA1_6 , \U4/DATA1_7 , \U4/DATA1_8 ,
         \U4/DATA1_9 , \U4/DATA1_10 , \U4/DATA1_11 , \U4/DATA1_12 ,
         \U4/DATA1_13 , \U4/DATA1_14 , \U4/DATA1_15 , \U4/DATA1_16 ,
         \U4/DATA1_17 , \U4/DATA1_18 , \U4/DATA1_19 , \U4/DATA1_20 ,
         \U4/DATA1_21 , \U4/DATA1_22 , \U4/DATA1_23 , \add_41/carry[4] ,
         \add_41/carry[3] , \add_41/carry[2] , \add_41/A[0] , \add_41/A[1] ,
         \add_41/A[2] , \add_41/A[3] , n1, n28, n32, n35, n41, n42, n43, n44,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n61, n65, n69,
         n73, n74, n75, n76, n77, n80, n84, n88, n92, n93, n96, n97, n100,
         n101, n104, n105, n108, n109, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n139,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n720, n721, n722, n723,
         n724, n725, n726, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814;
  assign \U12/DATA2_0  = Element[24];
  assign \U12/DATA2_1  = Element[25];
  assign \U12/DATA2_2  = Element[26];
  assign \U12/DATA2_3  = Element[27];
  assign \U12/DATA2_4  = Element[28];
  assign \U12/DATA2_5  = Element[29];
  assign \U12/DATA2_6  = Element[30];
  assign \U12/DATA2_7  = Element[31];
  assign \U12/DATA2_8  = Element[32];
  assign \U12/DATA2_9  = Element[33];
  assign \U12/DATA2_10  = Element[34];
  assign \U12/DATA2_11  = Element[35];
  assign \U12/DATA2_12  = Element[36];
  assign \U12/DATA2_13  = Element[37];
  assign \U12/DATA2_14  = Element[38];
  assign \U12/DATA2_15  = Element[39];
  assign \U12/DATA2_16  = Element[40];
  assign \U12/DATA2_17  = Element[41];
  assign \U12/DATA2_18  = Element[42];
  assign \U12/DATA2_19  = Element[43];
  assign \U12/DATA2_20  = Element[44];
  assign \U12/DATA2_21  = Element[45];
  assign \U12/DATA2_22  = Element[46];
  assign \U12/DATA2_23  = Element[47];
  assign \U12/DATA1_0  = Element[0];
  assign \U12/DATA1_1  = Element[1];
  assign \U12/DATA1_2  = Element[2];
  assign \U12/DATA1_3  = Element[3];
  assign \U12/DATA1_4  = Element[4];
  assign \U12/DATA1_5  = Element[5];
  assign \U12/DATA1_6  = Element[6];
  assign \U12/DATA1_7  = Element[7];
  assign \U12/DATA1_8  = Element[8];
  assign \U12/DATA1_9  = Element[9];
  assign \U12/DATA1_10  = Element[10];
  assign \U12/DATA1_11  = Element[11];
  assign \U12/DATA1_12  = Element[12];
  assign \U12/DATA1_13  = Element[13];
  assign \U12/DATA1_14  = Element[14];
  assign \U12/DATA1_15  = Element[15];
  assign \U12/DATA1_16  = Element[16];
  assign \U12/DATA1_17  = Element[17];
  assign \U12/DATA1_18  = Element[18];
  assign \U12/DATA1_19  = Element[19];
  assign \U12/DATA1_20  = Element[20];
  assign \U12/DATA1_21  = Element[21];
  assign \U12/DATA1_22  = Element[22];
  assign \U12/DATA1_23  = Element[23];
  assign \U11/DATA2_0  = NewElement[24];
  assign \U11/DATA2_1  = NewElement[25];
  assign \U11/DATA2_2  = NewElement[26];
  assign \U11/DATA2_3  = NewElement[27];
  assign \U11/DATA2_4  = NewElement[28];
  assign \U11/DATA2_5  = NewElement[29];
  assign \U11/DATA2_6  = NewElement[30];
  assign \U11/DATA2_7  = NewElement[31];
  assign \U11/DATA2_8  = NewElement[32];
  assign \U11/DATA2_9  = NewElement[33];
  assign \U11/DATA2_10  = NewElement[34];
  assign \U11/DATA2_11  = NewElement[35];
  assign \U11/DATA2_12  = NewElement[36];
  assign \U11/DATA2_13  = NewElement[37];
  assign \U11/DATA2_14  = NewElement[38];
  assign \U11/DATA2_15  = NewElement[39];
  assign \U11/DATA2_16  = NewElement[40];
  assign \U11/DATA2_17  = NewElement[41];
  assign \U11/DATA2_18  = NewElement[42];
  assign \U11/DATA2_19  = NewElement[43];
  assign \U11/DATA2_20  = NewElement[44];
  assign \U11/DATA2_21  = NewElement[45];
  assign \U11/DATA2_22  = NewElement[46];
  assign \U11/DATA2_23  = NewElement[47];
  assign \U11/DATA1_0  = NewElement[0];
  assign \U11/DATA1_1  = NewElement[1];
  assign \U11/DATA1_2  = NewElement[2];
  assign \U11/DATA1_3  = NewElement[3];
  assign \U11/DATA1_4  = NewElement[4];
  assign \U11/DATA1_5  = NewElement[5];
  assign \U11/DATA1_6  = NewElement[6];
  assign \U11/DATA1_7  = NewElement[7];
  assign \U11/DATA1_8  = NewElement[8];
  assign \U11/DATA1_9  = NewElement[9];
  assign \U11/DATA1_10  = NewElement[10];
  assign \U11/DATA1_11  = NewElement[11];
  assign \U11/DATA1_12  = NewElement[12];
  assign \U11/DATA1_13  = NewElement[13];
  assign \U11/DATA1_14  = NewElement[14];
  assign \U11/DATA1_15  = NewElement[15];
  assign \U11/DATA1_16  = NewElement[16];
  assign \U11/DATA1_17  = NewElement[17];
  assign \U11/DATA1_18  = NewElement[18];
  assign \U11/DATA1_19  = NewElement[19];
  assign \U11/DATA1_20  = NewElement[20];
  assign \U11/DATA1_21  = NewElement[21];
  assign \U11/DATA1_22  = NewElement[22];
  assign \U11/DATA1_23  = NewElement[23];
  assign SubInput1[0] = \U8/Z_0 ;
  assign SubInput1[1] = \U8/Z_1 ;
  assign SubInput1[2] = \U8/Z_2 ;
  assign SubInput1[3] = \U8/Z_3 ;
  assign SubInput1[4] = \U8/Z_4 ;
  assign SubInput1[5] = \U8/Z_5 ;
  assign SubInput1[6] = \U8/Z_6 ;
  assign SubInput1[7] = \U8/Z_7 ;
  assign SubInput1[8] = \U8/Z_8 ;
  assign SubInput1[9] = \U8/Z_9 ;
  assign SubInput1[10] = \U8/Z_10 ;
  assign SubInput1[11] = \U8/Z_11 ;
  assign SubInput1[12] = \U8/Z_12 ;
  assign SubInput1[13] = \U8/Z_13 ;
  assign SubInput1[14] = \U8/Z_14 ;
  assign SubInput1[15] = \U8/Z_15 ;
  assign SubInput1[16] = \U8/Z_16 ;
  assign SubInput1[17] = \U8/Z_17 ;
  assign SubInput1[18] = \U8/Z_18 ;
  assign SubInput1[19] = \U8/Z_19 ;
  assign SubInput1[20] = \U8/Z_20 ;
  assign SubInput1[21] = \U8/Z_21 ;
  assign SubInput1[22] = \U8/Z_22 ;
  assign SubInput1[23] = \U8/Z_23 ;
  assign SubInput2[0] = \U7/Z_0 ;
  assign SubInput2[1] = \U7/Z_1 ;
  assign SubInput2[2] = \U7/Z_2 ;
  assign SubInput2[3] = \U7/Z_3 ;
  assign SubInput2[4] = \U7/Z_4 ;
  assign SubInput2[5] = \U7/Z_5 ;
  assign SubInput2[6] = \U7/Z_6 ;
  assign SubInput2[7] = \U7/Z_7 ;
  assign SubInput2[8] = \U7/Z_8 ;
  assign SubInput2[9] = \U7/Z_9 ;
  assign SubInput2[10] = \U7/Z_10 ;
  assign SubInput2[11] = \U7/Z_11 ;
  assign SubInput2[12] = \U7/Z_12 ;
  assign SubInput2[13] = \U7/Z_13 ;
  assign SubInput2[14] = \U7/Z_14 ;
  assign SubInput2[15] = \U7/Z_15 ;
  assign SubInput2[16] = \U7/Z_16 ;
  assign SubInput2[17] = \U7/Z_17 ;
  assign SubInput2[18] = \U7/Z_18 ;
  assign SubInput2[19] = \U7/Z_19 ;
  assign SubInput2[20] = \U7/Z_20 ;
  assign SubInput2[21] = \U7/Z_21 ;
  assign SubInput2[22] = \U7/Z_22 ;
  assign SubInput2[23] = \U7/Z_23 ;
  assign \U6/DATA2_0  = DiagonalX[24];
  assign \U6/DATA2_1  = DiagonalX[25];
  assign \U6/DATA2_2  = DiagonalX[26];
  assign \U6/DATA2_3  = DiagonalX[27];
  assign \U6/DATA2_4  = DiagonalX[28];
  assign \U6/DATA2_5  = DiagonalX[29];
  assign \U6/DATA2_6  = DiagonalX[30];
  assign \U6/DATA2_7  = DiagonalX[31];
  assign \U6/DATA2_8  = DiagonalX[32];
  assign \U6/DATA2_9  = DiagonalX[33];
  assign \U6/DATA2_10  = DiagonalX[34];
  assign \U6/DATA2_11  = DiagonalX[35];
  assign \U6/DATA2_12  = DiagonalX[36];
  assign \U6/DATA2_13  = DiagonalX[37];
  assign \U6/DATA2_14  = DiagonalX[38];
  assign \U6/DATA2_15  = DiagonalX[39];
  assign \U6/DATA2_16  = DiagonalX[40];
  assign \U6/DATA2_17  = DiagonalX[41];
  assign \U6/DATA2_18  = DiagonalX[42];
  assign \U6/DATA2_19  = DiagonalX[43];
  assign \U6/DATA2_20  = DiagonalX[44];
  assign \U6/DATA2_21  = DiagonalX[45];
  assign \U6/DATA2_22  = DiagonalX[46];
  assign \U6/DATA2_23  = DiagonalX[47];
  assign \U6/DATA1_0  = DiagonalX[0];
  assign \U6/DATA1_1  = DiagonalX[1];
  assign \U6/DATA1_2  = DiagonalX[2];
  assign \U6/DATA1_3  = DiagonalX[3];
  assign \U6/DATA1_4  = DiagonalX[4];
  assign \U6/DATA1_5  = DiagonalX[5];
  assign \U6/DATA1_6  = DiagonalX[6];
  assign \U6/DATA1_7  = DiagonalX[7];
  assign \U6/DATA1_8  = DiagonalX[8];
  assign \U6/DATA1_9  = DiagonalX[9];
  assign \U6/DATA1_10  = DiagonalX[10];
  assign \U6/DATA1_11  = DiagonalX[11];
  assign \U6/DATA1_12  = DiagonalX[12];
  assign \U6/DATA1_13  = DiagonalX[13];
  assign \U6/DATA1_14  = DiagonalX[14];
  assign \U6/DATA1_15  = DiagonalX[15];
  assign \U6/DATA1_16  = DiagonalX[16];
  assign \U6/DATA1_17  = DiagonalX[17];
  assign \U6/DATA1_18  = DiagonalX[18];
  assign \U6/DATA1_19  = DiagonalX[19];
  assign \U6/DATA1_20  = DiagonalX[20];
  assign \U6/DATA1_21  = DiagonalX[21];
  assign \U6/DATA1_22  = DiagonalX[22];
  assign \U6/DATA1_23  = DiagonalX[23];
  assign \U5/DATA1_0  = DiagonalY[24];
  assign \U5/DATA1_1  = DiagonalY[25];
  assign \U5/DATA1_2  = DiagonalY[26];
  assign \U5/DATA1_3  = DiagonalY[27];
  assign \U5/DATA1_4  = DiagonalY[28];
  assign \U5/DATA1_5  = DiagonalY[29];
  assign \U5/DATA1_6  = DiagonalY[30];
  assign \U5/DATA1_7  = DiagonalY[31];
  assign \U5/DATA1_8  = DiagonalY[32];
  assign \U5/DATA1_9  = DiagonalY[33];
  assign \U5/DATA1_10  = DiagonalY[34];
  assign \U5/DATA1_11  = DiagonalY[35];
  assign \U5/DATA1_12  = DiagonalY[36];
  assign \U5/DATA1_13  = DiagonalY[37];
  assign \U5/DATA1_14  = DiagonalY[38];
  assign \U5/DATA1_15  = DiagonalY[39];
  assign \U5/DATA1_16  = DiagonalY[40];
  assign \U5/DATA1_17  = DiagonalY[41];
  assign \U5/DATA1_18  = DiagonalY[42];
  assign \U5/DATA1_19  = DiagonalY[43];
  assign \U5/DATA1_20  = DiagonalY[44];
  assign \U5/DATA1_21  = DiagonalY[45];
  assign \U5/DATA1_22  = DiagonalY[46];
  assign \U5/DATA1_23  = DiagonalY[47];
  assign AddInput1[0] = \U4/Z_0 ;
  assign AddInput1[1] = \U4/Z_1 ;
  assign AddInput1[2] = \U4/Z_2 ;
  assign AddInput1[3] = \U4/Z_3 ;
  assign AddInput1[4] = \U4/Z_4 ;
  assign AddInput1[5] = \U4/Z_5 ;
  assign AddInput1[6] = \U4/Z_6 ;
  assign AddInput1[7] = \U4/Z_7 ;
  assign AddInput1[8] = \U4/Z_8 ;
  assign AddInput1[9] = \U4/Z_9 ;
  assign AddInput1[10] = \U4/Z_10 ;
  assign AddInput1[11] = \U4/Z_11 ;
  assign AddInput1[12] = \U4/Z_12 ;
  assign AddInput1[13] = \U4/Z_13 ;
  assign AddInput1[14] = \U4/Z_14 ;
  assign AddInput1[15] = \U4/Z_15 ;
  assign AddInput1[16] = \U4/Z_16 ;
  assign AddInput1[17] = \U4/Z_17 ;
  assign AddInput1[18] = \U4/Z_18 ;
  assign AddInput1[19] = \U4/Z_19 ;
  assign AddInput1[20] = \U4/Z_20 ;
  assign AddInput1[21] = \U4/Z_21 ;
  assign AddInput1[22] = \U4/Z_22 ;
  assign AddInput1[23] = \U4/Z_23 ;
  assign \U4/DATA1_0  = DiagonalY[0];
  assign \U4/DATA1_1  = DiagonalY[1];
  assign \U4/DATA1_2  = DiagonalY[2];
  assign \U4/DATA1_3  = DiagonalY[3];
  assign \U4/DATA1_4  = DiagonalY[4];
  assign \U4/DATA1_5  = DiagonalY[5];
  assign \U4/DATA1_6  = DiagonalY[6];
  assign \U4/DATA1_7  = DiagonalY[7];
  assign \U4/DATA1_8  = DiagonalY[8];
  assign \U4/DATA1_9  = DiagonalY[9];
  assign \U4/DATA1_10  = DiagonalY[10];
  assign \U4/DATA1_11  = DiagonalY[11];
  assign \U4/DATA1_12  = DiagonalY[12];
  assign \U4/DATA1_13  = DiagonalY[13];
  assign \U4/DATA1_14  = DiagonalY[14];
  assign \U4/DATA1_15  = DiagonalY[15];
  assign \U4/DATA1_16  = DiagonalY[16];
  assign \U4/DATA1_17  = DiagonalY[17];
  assign \U4/DATA1_18  = DiagonalY[18];
  assign \U4/DATA1_19  = DiagonalY[19];
  assign \U4/DATA1_20  = DiagonalY[20];
  assign \U4/DATA1_21  = DiagonalY[21];
  assign \U4/DATA1_22  = DiagonalY[22];
  assign \U4/DATA1_23  = DiagonalY[23];

  HA_X1 \add_41/U1_1_1  ( .A(\add_41/A[1] ), .B(\add_41/A[0] ), .CO(
        \add_41/carry[2] ), .S(\U3/U1/DATA2_1 ) );
  HA_X1 \add_41/U1_1_2  ( .A(\add_41/A[2] ), .B(\add_41/carry[2] ), .CO(
        \add_41/carry[3] ), .S(\U3/U1/DATA2_2 ) );
  HA_X1 \add_41/U1_1_3  ( .A(\add_41/A[3] ), .B(\add_41/carry[3] ), .CO(
        \add_41/carry[4] ), .S(\U3/U1/DATA2_3 ) );
  DFF_X1 \Count_reg[0]  ( .D(n757), .CK(clock), .Q(\add_41/A[0] ), .QN(n386)
         );
  DFF_X1 \Count_reg[1]  ( .D(n390), .CK(clock), .Q(\add_41/A[1] ), .QN(n385)
         );
  DFF_X1 \Count_reg[2]  ( .D(n389), .CK(clock), .Q(\add_41/A[2] ), .QN(n384)
         );
  DFF_X1 \Count_reg[3]  ( .D(n388), .CK(clock), .Q(\add_41/A[3] ), .QN(n383)
         );
  DFF_X1 \NewDiagonalX_reg[47]  ( .D(n380), .CK(clock), .Q(NewDiagonalX[47]), 
        .QN(n284) );
  DFF_X1 \NewDiagonalX_reg[46]  ( .D(n379), .CK(clock), .Q(NewDiagonalX[46]), 
        .QN(n283) );
  DFF_X1 \NewDiagonalX_reg[45]  ( .D(n378), .CK(clock), .Q(NewDiagonalX[45]), 
        .QN(n282) );
  DFF_X1 \NewDiagonalX_reg[44]  ( .D(n377), .CK(clock), .Q(NewDiagonalX[44]), 
        .QN(n281) );
  DFF_X1 \NewDiagonalX_reg[43]  ( .D(n376), .CK(clock), .Q(NewDiagonalX[43]), 
        .QN(n280) );
  DFF_X1 \NewDiagonalX_reg[42]  ( .D(n375), .CK(clock), .Q(NewDiagonalX[42]), 
        .QN(n279) );
  DFF_X1 \NewDiagonalX_reg[41]  ( .D(n374), .CK(clock), .Q(NewDiagonalX[41]), 
        .QN(n278) );
  DFF_X1 \NewDiagonalX_reg[40]  ( .D(n373), .CK(clock), .Q(NewDiagonalX[40]), 
        .QN(n277) );
  DFF_X1 \NewDiagonalX_reg[39]  ( .D(n372), .CK(clock), .Q(NewDiagonalX[39]), 
        .QN(n276) );
  DFF_X1 \NewDiagonalX_reg[38]  ( .D(n371), .CK(clock), .Q(NewDiagonalX[38]), 
        .QN(n275) );
  DFF_X1 \NewDiagonalX_reg[37]  ( .D(n370), .CK(clock), .Q(NewDiagonalX[37]), 
        .QN(n274) );
  DFF_X1 \NewDiagonalX_reg[36]  ( .D(n369), .CK(clock), .Q(NewDiagonalX[36]), 
        .QN(n273) );
  DFF_X1 \NewDiagonalX_reg[35]  ( .D(n368), .CK(clock), .Q(NewDiagonalX[35]), 
        .QN(n272) );
  DFF_X1 \NewDiagonalX_reg[34]  ( .D(n367), .CK(clock), .Q(NewDiagonalX[34]), 
        .QN(n271) );
  DFF_X1 \NewDiagonalX_reg[33]  ( .D(n366), .CK(clock), .Q(NewDiagonalX[33]), 
        .QN(n270) );
  DFF_X1 \NewDiagonalX_reg[32]  ( .D(n365), .CK(clock), .Q(NewDiagonalX[32]), 
        .QN(n269) );
  DFF_X1 \NewDiagonalX_reg[31]  ( .D(n364), .CK(clock), .Q(NewDiagonalX[31]), 
        .QN(n268) );
  DFF_X1 \NewDiagonalX_reg[30]  ( .D(n363), .CK(clock), .Q(NewDiagonalX[30]), 
        .QN(n267) );
  DFF_X1 \NewDiagonalX_reg[29]  ( .D(n362), .CK(clock), .Q(NewDiagonalX[29]), 
        .QN(n266) );
  DFF_X1 \NewDiagonalX_reg[28]  ( .D(n361), .CK(clock), .Q(NewDiagonalX[28]), 
        .QN(n265) );
  DFF_X1 \NewDiagonalX_reg[27]  ( .D(n360), .CK(clock), .Q(NewDiagonalX[27]), 
        .QN(n264) );
  DFF_X1 \NewDiagonalX_reg[26]  ( .D(n359), .CK(clock), .Q(NewDiagonalX[26]), 
        .QN(n263) );
  DFF_X1 \NewDiagonalX_reg[25]  ( .D(n358), .CK(clock), .Q(NewDiagonalX[25]), 
        .QN(n262) );
  DFF_X1 \NewDiagonalX_reg[24]  ( .D(n357), .CK(clock), .Q(NewDiagonalX[24]), 
        .QN(n261) );
  DFF_X1 \NewDiagonalY_reg[47]  ( .D(n356), .CK(clock), .Q(NewDiagonalY[47]), 
        .QN(n260) );
  DFF_X1 \NewDiagonalY_reg[46]  ( .D(n355), .CK(clock), .Q(NewDiagonalY[46]), 
        .QN(n259) );
  DFF_X1 \NewDiagonalY_reg[45]  ( .D(n354), .CK(clock), .Q(NewDiagonalY[45]), 
        .QN(n258) );
  DFF_X1 \NewDiagonalY_reg[44]  ( .D(n353), .CK(clock), .Q(NewDiagonalY[44]), 
        .QN(n257) );
  DFF_X1 \NewDiagonalY_reg[43]  ( .D(n352), .CK(clock), .Q(NewDiagonalY[43]), 
        .QN(n256) );
  DFF_X1 \NewDiagonalY_reg[42]  ( .D(n351), .CK(clock), .Q(NewDiagonalY[42]), 
        .QN(n255) );
  DFF_X1 \NewDiagonalY_reg[41]  ( .D(n350), .CK(clock), .Q(NewDiagonalY[41]), 
        .QN(n254) );
  DFF_X1 \NewDiagonalY_reg[40]  ( .D(n349), .CK(clock), .Q(NewDiagonalY[40]), 
        .QN(n253) );
  DFF_X1 \NewDiagonalY_reg[39]  ( .D(n348), .CK(clock), .Q(NewDiagonalY[39]), 
        .QN(n252) );
  DFF_X1 \NewDiagonalY_reg[38]  ( .D(n347), .CK(clock), .Q(NewDiagonalY[38]), 
        .QN(n251) );
  DFF_X1 \NewDiagonalY_reg[37]  ( .D(n346), .CK(clock), .Q(NewDiagonalY[37]), 
        .QN(n250) );
  DFF_X1 \NewDiagonalY_reg[36]  ( .D(n345), .CK(clock), .Q(NewDiagonalY[36]), 
        .QN(n249) );
  DFF_X1 \NewDiagonalY_reg[35]  ( .D(n344), .CK(clock), .Q(NewDiagonalY[35]), 
        .QN(n248) );
  DFF_X1 \NewDiagonalY_reg[34]  ( .D(n343), .CK(clock), .Q(NewDiagonalY[34]), 
        .QN(n247) );
  DFF_X1 \NewDiagonalY_reg[33]  ( .D(n342), .CK(clock), .Q(NewDiagonalY[33]), 
        .QN(n246) );
  DFF_X1 \NewDiagonalY_reg[32]  ( .D(n341), .CK(clock), .Q(NewDiagonalY[32]), 
        .QN(n245) );
  DFF_X1 \NewDiagonalY_reg[31]  ( .D(n340), .CK(clock), .Q(NewDiagonalY[31]), 
        .QN(n244) );
  DFF_X1 \NewDiagonalY_reg[30]  ( .D(n339), .CK(clock), .Q(NewDiagonalY[30]), 
        .QN(n243) );
  DFF_X1 \NewDiagonalY_reg[29]  ( .D(n338), .CK(clock), .Q(NewDiagonalY[29]), 
        .QN(n242) );
  DFF_X1 \NewDiagonalY_reg[28]  ( .D(n337), .CK(clock), .Q(NewDiagonalY[28]), 
        .QN(n241) );
  DFF_X1 \NewDiagonalY_reg[27]  ( .D(n336), .CK(clock), .Q(NewDiagonalY[27]), 
        .QN(n240) );
  DFF_X1 \NewDiagonalY_reg[26]  ( .D(n335), .CK(clock), .Q(NewDiagonalY[26]), 
        .QN(n239) );
  DFF_X1 \NewDiagonalY_reg[25]  ( .D(n334), .CK(clock), .Q(NewDiagonalY[25]), 
        .QN(n238) );
  DFF_X1 \NewDiagonalY_reg[24]  ( .D(n333), .CK(clock), .Q(NewDiagonalY[24]), 
        .QN(n237) );
  DFF_X1 \NewDiagonalY_reg[23]  ( .D(n332), .CK(clock), .Q(NewDiagonalY[23]), 
        .QN(n236) );
  DFF_X1 \NewDiagonalY_reg[22]  ( .D(n331), .CK(clock), .Q(NewDiagonalY[22]), 
        .QN(n235) );
  DFF_X1 \NewDiagonalY_reg[21]  ( .D(n330), .CK(clock), .Q(NewDiagonalY[21]), 
        .QN(n234) );
  DFF_X1 \NewDiagonalY_reg[20]  ( .D(n329), .CK(clock), .Q(NewDiagonalY[20]), 
        .QN(n233) );
  DFF_X1 \NewDiagonalY_reg[19]  ( .D(n328), .CK(clock), .Q(NewDiagonalY[19]), 
        .QN(n232) );
  DFF_X1 \NewDiagonalY_reg[18]  ( .D(n327), .CK(clock), .Q(NewDiagonalY[18]), 
        .QN(n231) );
  DFF_X1 \NewDiagonalY_reg[17]  ( .D(n326), .CK(clock), .Q(NewDiagonalY[17]), 
        .QN(n230) );
  DFF_X1 \NewDiagonalY_reg[16]  ( .D(n325), .CK(clock), .Q(NewDiagonalY[16]), 
        .QN(n229) );
  DFF_X1 \NewDiagonalY_reg[15]  ( .D(n324), .CK(clock), .Q(NewDiagonalY[15]), 
        .QN(n228) );
  DFF_X1 \NewDiagonalY_reg[14]  ( .D(n323), .CK(clock), .Q(NewDiagonalY[14]), 
        .QN(n227) );
  DFF_X1 \NewDiagonalY_reg[13]  ( .D(n322), .CK(clock), .Q(NewDiagonalY[13]), 
        .QN(n226) );
  DFF_X1 \NewDiagonalY_reg[12]  ( .D(n321), .CK(clock), .Q(NewDiagonalY[12]), 
        .QN(n225) );
  DFF_X1 \NewDiagonalY_reg[11]  ( .D(n320), .CK(clock), .Q(NewDiagonalY[11]), 
        .QN(n224) );
  DFF_X1 \NewDiagonalY_reg[10]  ( .D(n319), .CK(clock), .Q(NewDiagonalY[10]), 
        .QN(n223) );
  DFF_X1 \NewDiagonalY_reg[9]  ( .D(n318), .CK(clock), .Q(NewDiagonalY[9]), 
        .QN(n222) );
  DFF_X1 \NewDiagonalY_reg[8]  ( .D(n317), .CK(clock), .Q(NewDiagonalY[8]), 
        .QN(n221) );
  DFF_X1 \NewDiagonalY_reg[7]  ( .D(n316), .CK(clock), .Q(NewDiagonalY[7]), 
        .QN(n220) );
  DFF_X1 \NewDiagonalY_reg[6]  ( .D(n315), .CK(clock), .Q(NewDiagonalY[6]), 
        .QN(n219) );
  DFF_X1 \NewDiagonalY_reg[5]  ( .D(n314), .CK(clock), .Q(NewDiagonalY[5]), 
        .QN(n218) );
  DFF_X1 \NewDiagonalY_reg[4]  ( .D(n313), .CK(clock), .Q(NewDiagonalY[4]), 
        .QN(n217) );
  DFF_X1 \NewDiagonalY_reg[3]  ( .D(n312), .CK(clock), .Q(NewDiagonalY[3]), 
        .QN(n216) );
  DFF_X1 \NewDiagonalY_reg[2]  ( .D(n311), .CK(clock), .Q(NewDiagonalY[2]), 
        .QN(n215) );
  DFF_X1 \NewDiagonalY_reg[1]  ( .D(n310), .CK(clock), .Q(NewDiagonalY[1]), 
        .QN(n214) );
  DFF_X1 \NewDiagonalY_reg[0]  ( .D(n309), .CK(clock), .Q(NewDiagonalY[0]), 
        .QN(n213) );
  DFF_X1 \NewDiagonalX_reg[23]  ( .D(n308), .CK(clock), .Q(NewDiagonalX[23]), 
        .QN(n212) );
  DFF_X1 \NewDiagonalX_reg[22]  ( .D(n307), .CK(clock), .Q(NewDiagonalX[22]), 
        .QN(n211) );
  DFF_X1 \NewDiagonalX_reg[21]  ( .D(n306), .CK(clock), .Q(NewDiagonalX[21]), 
        .QN(n210) );
  DFF_X1 \NewDiagonalX_reg[20]  ( .D(n305), .CK(clock), .Q(NewDiagonalX[20]), 
        .QN(n209) );
  DFF_X1 \NewDiagonalX_reg[19]  ( .D(n304), .CK(clock), .Q(NewDiagonalX[19]), 
        .QN(n208) );
  DFF_X1 \NewDiagonalX_reg[18]  ( .D(n303), .CK(clock), .Q(NewDiagonalX[18]), 
        .QN(n207) );
  DFF_X1 \NewDiagonalX_reg[17]  ( .D(n302), .CK(clock), .Q(NewDiagonalX[17]), 
        .QN(n206) );
  DFF_X1 \NewDiagonalX_reg[16]  ( .D(n301), .CK(clock), .Q(NewDiagonalX[16]), 
        .QN(n205) );
  DFF_X1 \NewDiagonalX_reg[15]  ( .D(n300), .CK(clock), .Q(NewDiagonalX[15]), 
        .QN(n204) );
  DFF_X1 \NewDiagonalX_reg[14]  ( .D(n299), .CK(clock), .Q(NewDiagonalX[14]), 
        .QN(n203) );
  DFF_X1 \NewDiagonalX_reg[13]  ( .D(n298), .CK(clock), .Q(NewDiagonalX[13]), 
        .QN(n202) );
  DFF_X1 \NewDiagonalX_reg[12]  ( .D(n297), .CK(clock), .Q(NewDiagonalX[12]), 
        .QN(n201) );
  DFF_X1 \NewDiagonalX_reg[11]  ( .D(n296), .CK(clock), .Q(NewDiagonalX[11]), 
        .QN(n200) );
  DFF_X1 \NewDiagonalX_reg[10]  ( .D(n295), .CK(clock), .Q(NewDiagonalX[10]), 
        .QN(n199) );
  DFF_X1 \NewDiagonalX_reg[9]  ( .D(n294), .CK(clock), .Q(NewDiagonalX[9]), 
        .QN(n198) );
  DFF_X1 \NewDiagonalX_reg[8]  ( .D(n293), .CK(clock), .Q(NewDiagonalX[8]), 
        .QN(n197) );
  DFF_X1 \NewDiagonalX_reg[7]  ( .D(n292), .CK(clock), .Q(NewDiagonalX[7]), 
        .QN(n196) );
  DFF_X1 \NewDiagonalX_reg[6]  ( .D(n291), .CK(clock), .Q(NewDiagonalX[6]), 
        .QN(n195) );
  DFF_X1 \NewDiagonalX_reg[5]  ( .D(n290), .CK(clock), .Q(NewDiagonalX[5]), 
        .QN(n194) );
  DFF_X1 \NewDiagonalX_reg[4]  ( .D(n289), .CK(clock), .Q(NewDiagonalX[4]), 
        .QN(n193) );
  DFF_X1 \NewDiagonalX_reg[3]  ( .D(n288), .CK(clock), .Q(NewDiagonalX[3]), 
        .QN(n192) );
  DFF_X1 \NewDiagonalX_reg[2]  ( .D(n287), .CK(clock), .Q(NewDiagonalX[2]), 
        .QN(n191) );
  DFF_X1 \NewDiagonalX_reg[1]  ( .D(n286), .CK(clock), .Q(NewDiagonalX[1]), 
        .QN(n190) );
  DFF_X1 \NewDiagonalX_reg[0]  ( .D(n285), .CK(clock), .Q(NewDiagonalX[0]), 
        .QN(n189) );
  DFF_X1 DiagonalXDone_reg ( .D(n381), .CK(clock), .Q(DiagonalXDone), .QN(n720) );
  OAI22_X2 U3 ( .A1(n1), .A2(n814), .B1(n189), .B2(n756), .ZN(n285) );
  OAI22_X2 U4 ( .A1(n1), .A2(n813), .B1(n190), .B2(n756), .ZN(n286) );
  OAI22_X2 U5 ( .A1(n1), .A2(n812), .B1(n191), .B2(n756), .ZN(n287) );
  OAI22_X2 U6 ( .A1(n1), .A2(n811), .B1(n192), .B2(n756), .ZN(n288) );
  OAI22_X2 U7 ( .A1(n1), .A2(n810), .B1(n193), .B2(n756), .ZN(n289) );
  OAI22_X2 U8 ( .A1(n1), .A2(n809), .B1(n194), .B2(n756), .ZN(n290) );
  OAI22_X2 U9 ( .A1(n1), .A2(n808), .B1(n195), .B2(n756), .ZN(n291) );
  OAI22_X2 U10 ( .A1(n1), .A2(n807), .B1(n196), .B2(n756), .ZN(n292) );
  OAI22_X2 U11 ( .A1(n1), .A2(n806), .B1(n197), .B2(n756), .ZN(n293) );
  OAI22_X2 U12 ( .A1(n1), .A2(n805), .B1(n198), .B2(n756), .ZN(n294) );
  OAI22_X2 U13 ( .A1(n1), .A2(n804), .B1(n199), .B2(n756), .ZN(n295) );
  OAI22_X2 U14 ( .A1(n1), .A2(n803), .B1(n200), .B2(n756), .ZN(n296) );
  OAI22_X2 U15 ( .A1(n1), .A2(n802), .B1(n201), .B2(n756), .ZN(n297) );
  OAI22_X2 U16 ( .A1(n1), .A2(n801), .B1(n202), .B2(n756), .ZN(n298) );
  OAI22_X2 U17 ( .A1(n1), .A2(n800), .B1(n203), .B2(n756), .ZN(n299) );
  OAI22_X2 U18 ( .A1(n1), .A2(n799), .B1(n204), .B2(n756), .ZN(n300) );
  OAI22_X2 U19 ( .A1(n1), .A2(n798), .B1(n205), .B2(n756), .ZN(n301) );
  OAI22_X2 U20 ( .A1(n1), .A2(n797), .B1(n206), .B2(n756), .ZN(n302) );
  OAI22_X2 U21 ( .A1(n1), .A2(n796), .B1(n207), .B2(n756), .ZN(n303) );
  OAI22_X2 U22 ( .A1(n1), .A2(n795), .B1(n208), .B2(n756), .ZN(n304) );
  OAI22_X2 U23 ( .A1(n1), .A2(n794), .B1(n209), .B2(n756), .ZN(n305) );
  OAI22_X2 U24 ( .A1(n1), .A2(n793), .B1(n210), .B2(n756), .ZN(n306) );
  OAI22_X2 U25 ( .A1(n1), .A2(n792), .B1(n211), .B2(n756), .ZN(n307) );
  OAI22_X2 U26 ( .A1(n1), .A2(n791), .B1(n212), .B2(n756), .ZN(n308) );
  OAI22_X2 U28 ( .A1(n814), .A2(n755), .B1(n213), .B2(n28), .ZN(n309) );
  OAI22_X2 U29 ( .A1(n813), .A2(n755), .B1(n214), .B2(n28), .ZN(n310) );
  OAI22_X2 U30 ( .A1(n812), .A2(n755), .B1(n215), .B2(n28), .ZN(n311) );
  OAI22_X2 U31 ( .A1(n811), .A2(n755), .B1(n216), .B2(n28), .ZN(n312) );
  OAI22_X2 U32 ( .A1(n810), .A2(n755), .B1(n217), .B2(n28), .ZN(n313) );
  OAI22_X2 U33 ( .A1(n809), .A2(n755), .B1(n218), .B2(n28), .ZN(n314) );
  OAI22_X2 U34 ( .A1(n808), .A2(n755), .B1(n219), .B2(n28), .ZN(n315) );
  OAI22_X2 U35 ( .A1(n807), .A2(n755), .B1(n220), .B2(n28), .ZN(n316) );
  OAI22_X2 U36 ( .A1(n806), .A2(n755), .B1(n221), .B2(n754), .ZN(n317) );
  OAI22_X2 U37 ( .A1(n805), .A2(n755), .B1(n222), .B2(n754), .ZN(n318) );
  OAI22_X2 U38 ( .A1(n804), .A2(n755), .B1(n223), .B2(n754), .ZN(n319) );
  OAI22_X2 U39 ( .A1(n803), .A2(n755), .B1(n224), .B2(n754), .ZN(n320) );
  OAI22_X2 U40 ( .A1(n802), .A2(n755), .B1(n225), .B2(n754), .ZN(n321) );
  OAI22_X2 U41 ( .A1(n801), .A2(n755), .B1(n226), .B2(n754), .ZN(n322) );
  OAI22_X2 U42 ( .A1(n800), .A2(n755), .B1(n227), .B2(n754), .ZN(n323) );
  OAI22_X2 U43 ( .A1(n799), .A2(n755), .B1(n228), .B2(n754), .ZN(n324) );
  OAI22_X2 U44 ( .A1(n798), .A2(n755), .B1(n229), .B2(n754), .ZN(n325) );
  OAI22_X2 U45 ( .A1(n797), .A2(n755), .B1(n230), .B2(n754), .ZN(n326) );
  OAI22_X2 U46 ( .A1(n796), .A2(n755), .B1(n231), .B2(n754), .ZN(n327) );
  OAI22_X2 U47 ( .A1(n795), .A2(n755), .B1(n232), .B2(n754), .ZN(n328) );
  OAI22_X2 U48 ( .A1(n794), .A2(n755), .B1(n233), .B2(n754), .ZN(n329) );
  OAI22_X2 U49 ( .A1(n793), .A2(n755), .B1(n234), .B2(n754), .ZN(n330) );
  OAI22_X2 U50 ( .A1(n792), .A2(n755), .B1(n235), .B2(n754), .ZN(n331) );
  OAI22_X2 U51 ( .A1(n791), .A2(n755), .B1(n236), .B2(n754), .ZN(n332) );
  OAI22_X2 U55 ( .A1(n814), .A2(n753), .B1(n237), .B2(n723), .ZN(n333) );
  OAI22_X2 U56 ( .A1(n813), .A2(n753), .B1(n238), .B2(n723), .ZN(n334) );
  OAI22_X2 U57 ( .A1(n812), .A2(n753), .B1(n239), .B2(n723), .ZN(n335) );
  OAI22_X2 U58 ( .A1(n811), .A2(n753), .B1(n240), .B2(n723), .ZN(n336) );
  OAI22_X2 U59 ( .A1(n810), .A2(n753), .B1(n241), .B2(n723), .ZN(n337) );
  OAI22_X2 U60 ( .A1(n809), .A2(n753), .B1(n242), .B2(n723), .ZN(n338) );
  OAI22_X2 U61 ( .A1(n808), .A2(n753), .B1(n243), .B2(n723), .ZN(n339) );
  OAI22_X2 U62 ( .A1(n807), .A2(n753), .B1(n244), .B2(n723), .ZN(n340) );
  OAI22_X2 U63 ( .A1(n806), .A2(n753), .B1(n245), .B2(n723), .ZN(n341) );
  OAI22_X2 U64 ( .A1(n805), .A2(n753), .B1(n246), .B2(n723), .ZN(n342) );
  OAI22_X2 U65 ( .A1(n804), .A2(n753), .B1(n247), .B2(n723), .ZN(n343) );
  OAI22_X2 U66 ( .A1(n803), .A2(n753), .B1(n248), .B2(n723), .ZN(n344) );
  OAI22_X2 U67 ( .A1(n802), .A2(n753), .B1(n249), .B2(n723), .ZN(n345) );
  OAI22_X2 U68 ( .A1(n801), .A2(n753), .B1(n250), .B2(n723), .ZN(n346) );
  OAI22_X2 U69 ( .A1(n800), .A2(n753), .B1(n251), .B2(n723), .ZN(n347) );
  OAI22_X2 U70 ( .A1(n799), .A2(n753), .B1(n252), .B2(n723), .ZN(n348) );
  OAI22_X2 U71 ( .A1(n798), .A2(n753), .B1(n253), .B2(n723), .ZN(n349) );
  OAI22_X2 U72 ( .A1(n797), .A2(n753), .B1(n254), .B2(n723), .ZN(n350) );
  OAI22_X2 U73 ( .A1(n796), .A2(n753), .B1(n255), .B2(n723), .ZN(n351) );
  OAI22_X2 U74 ( .A1(n795), .A2(n753), .B1(n256), .B2(n723), .ZN(n352) );
  OAI22_X2 U75 ( .A1(n794), .A2(n753), .B1(n257), .B2(n723), .ZN(n353) );
  OAI22_X2 U76 ( .A1(n793), .A2(n753), .B1(n258), .B2(n723), .ZN(n354) );
  OAI22_X2 U77 ( .A1(n792), .A2(n753), .B1(n259), .B2(n723), .ZN(n355) );
  OAI22_X2 U78 ( .A1(n791), .A2(n753), .B1(n260), .B2(n723), .ZN(n356) );
  OAI22_X2 U81 ( .A1(n814), .A2(n752), .B1(n261), .B2(n725), .ZN(n357) );
  OAI22_X2 U83 ( .A1(n813), .A2(n752), .B1(n262), .B2(n725), .ZN(n358) );
  OAI22_X2 U85 ( .A1(n812), .A2(n752), .B1(n263), .B2(n725), .ZN(n359) );
  OAI22_X2 U87 ( .A1(n811), .A2(n752), .B1(n264), .B2(n725), .ZN(n360) );
  OAI22_X2 U89 ( .A1(n810), .A2(n752), .B1(n265), .B2(n725), .ZN(n361) );
  OAI22_X2 U91 ( .A1(n809), .A2(n752), .B1(n266), .B2(n725), .ZN(n362) );
  OAI22_X2 U93 ( .A1(n808), .A2(n752), .B1(n267), .B2(n725), .ZN(n363) );
  OAI22_X2 U95 ( .A1(n807), .A2(n752), .B1(n268), .B2(n725), .ZN(n364) );
  OAI22_X2 U97 ( .A1(n806), .A2(n752), .B1(n269), .B2(n725), .ZN(n365) );
  OAI22_X2 U99 ( .A1(n805), .A2(n752), .B1(n270), .B2(n725), .ZN(n366) );
  OAI22_X2 U101 ( .A1(n804), .A2(n752), .B1(n271), .B2(n725), .ZN(n367) );
  OAI22_X2 U103 ( .A1(n803), .A2(n752), .B1(n272), .B2(n725), .ZN(n368) );
  OAI22_X2 U105 ( .A1(n802), .A2(n752), .B1(n273), .B2(n725), .ZN(n369) );
  OAI22_X2 U107 ( .A1(n801), .A2(n752), .B1(n274), .B2(n725), .ZN(n370) );
  OAI22_X2 U109 ( .A1(n800), .A2(n752), .B1(n275), .B2(n725), .ZN(n371) );
  OAI22_X2 U111 ( .A1(n799), .A2(n752), .B1(n276), .B2(n725), .ZN(n372) );
  OAI22_X2 U113 ( .A1(n798), .A2(n752), .B1(n277), .B2(n725), .ZN(n373) );
  OAI22_X2 U115 ( .A1(n797), .A2(n752), .B1(n278), .B2(n725), .ZN(n374) );
  OAI22_X2 U117 ( .A1(n796), .A2(n752), .B1(n279), .B2(n725), .ZN(n375) );
  OAI22_X2 U119 ( .A1(n795), .A2(n752), .B1(n280), .B2(n725), .ZN(n376) );
  OAI22_X2 U121 ( .A1(n794), .A2(n752), .B1(n281), .B2(n725), .ZN(n377) );
  OAI22_X2 U123 ( .A1(n793), .A2(n752), .B1(n282), .B2(n725), .ZN(n378) );
  OAI22_X2 U125 ( .A1(n792), .A2(n752), .B1(n283), .B2(n725), .ZN(n379) );
  OAI22_X2 U127 ( .A1(n791), .A2(n752), .B1(n284), .B2(n725), .ZN(n380) );
  NAND3_X2 U134 ( .A1(n35), .A2(\add_41/A[1] ), .A3(n386), .ZN(n1) );
  NAND2_X2 U135 ( .A1(n41), .A2(n42), .ZN(n387) );
  NAND3_X2 U136 ( .A1(n43), .A2(n382), .A3(\add_41/carry[4] ), .ZN(n42) );
  NOR3_X2 U138 ( .A1(EnableChange), .A2(reset), .A3(\add_41/carry[4] ), .ZN(
        n44) );
  NAND2_X2 U140 ( .A1(\U3/U1/DATA2_3 ), .A2(n43), .ZN(n48) );
  NAND2_X2 U142 ( .A1(\U3/U1/DATA2_2 ), .A2(n43), .ZN(n49) );
  NAND2_X2 U144 ( .A1(\U3/U1/DATA2_1 ), .A2(n43), .ZN(n50) );
  NOR3_X2 U147 ( .A1(EnableChange), .A2(reset), .A3(n759), .ZN(n43) );
  NAND2_X2 U149 ( .A1(n52), .A2(n53), .ZN(n47) );
  NOR4_X2 U150 ( .A1(n54), .A2(n55), .A3(n56), .A4(n57), .ZN(n53) );
  NAND4_X2 U151 ( .A1(n773), .A2(n767), .A3(n774), .A4(n61), .ZN(n57) );
  NOR3_X2 U152 ( .A1(\U12/DATA2_11 ), .A2(\U12/DATA2_13 ), .A3(\U12/DATA2_12 ), 
        .ZN(n61) );
  NAND4_X2 U153 ( .A1(n764), .A2(n763), .A3(n765), .A4(n65), .ZN(n56) );
  NOR3_X2 U154 ( .A1(\U12/DATA2_17 ), .A2(\U12/DATA2_19 ), .A3(\U12/DATA2_18 ), 
        .ZN(n65) );
  NAND4_X2 U155 ( .A1(n761), .A2(n760), .A3(n772), .A4(n69), .ZN(n55) );
  NOR3_X2 U156 ( .A1(\U12/DATA2_22 ), .A2(\U12/DATA2_3 ), .A3(\U12/DATA2_23 ), 
        .ZN(n69) );
  NAND4_X2 U157 ( .A1(n769), .A2(n768), .A3(n770), .A4(n73), .ZN(n54) );
  NOR4_X2 U158 ( .A1(reset), .A2(\U12/DATA2_9 ), .A3(\U12/DATA2_8 ), .A4(
        \U12/DATA2_7 ), .ZN(n73) );
  NOR4_X2 U159 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(n52) );
  NAND4_X2 U160 ( .A1(n789), .A2(n788), .A3(n790), .A4(n80), .ZN(n77) );
  NOR3_X2 U161 ( .A1(\U12/DATA1_10 ), .A2(\U12/DATA1_12 ), .A3(\U12/DATA1_11 ), 
        .ZN(n80) );
  NAND4_X2 U163 ( .A1(n780), .A2(n779), .A3(n781), .A4(n84), .ZN(n76) );
  NOR3_X2 U164 ( .A1(\U12/DATA1_16 ), .A2(\U12/DATA1_18 ), .A3(\U12/DATA1_17 ), 
        .ZN(n84) );
  NAND4_X2 U165 ( .A1(n787), .A2(n776), .A3(n777), .A4(n88), .ZN(n75) );
  NOR3_X2 U166 ( .A1(\U12/DATA1_21 ), .A2(\U12/DATA1_23 ), .A3(\U12/DATA1_22 ), 
        .ZN(n88) );
  NAND4_X2 U167 ( .A1(n785), .A2(n784), .A3(n786), .A4(n92), .ZN(n74) );
  NOR4_X2 U168 ( .A1(\U12/DATA1_9 ), .A2(\U12/DATA1_8 ), .A3(\U12/DATA1_7 ), 
        .A4(\U12/DATA1_6 ), .ZN(n92) );
  INV_X4 U169 ( .A(n93), .ZN(\U8/Z_9 ) );
  INV_X4 U171 ( .A(n96), .ZN(\U8/Z_8 ) );
  INV_X4 U173 ( .A(n97), .ZN(\U8/Z_7 ) );
  OAI22_X2 U175 ( .A1(n724), .A2(n768), .B1(n751), .B2(n783), .ZN(\U8/Z_6 ) );
  OAI22_X2 U178 ( .A1(n724), .A2(n769), .B1(n751), .B2(n784), .ZN(\U8/Z_5 ) );
  OAI22_X2 U181 ( .A1(n724), .A2(n770), .B1(n751), .B2(n785), .ZN(\U8/Z_4 ) );
  OAI22_X2 U184 ( .A1(n724), .A2(n771), .B1(n751), .B2(n786), .ZN(\U8/Z_3 ) );
  INV_X4 U187 ( .A(n100), .ZN(\U8/Z_23 ) );
  INV_X4 U189 ( .A(n101), .ZN(\U8/Z_22 ) );
  OAI22_X2 U191 ( .A1(n724), .A2(n760), .B1(n751), .B2(n775), .ZN(\U8/Z_21 )
         );
  OAI22_X2 U194 ( .A1(n724), .A2(n761), .B1(n751), .B2(n776), .ZN(\U8/Z_20 )
         );
  OAI22_X2 U197 ( .A1(n724), .A2(n772), .B1(n751), .B2(n787), .ZN(\U8/Z_2 ) );
  OAI22_X2 U200 ( .A1(n724), .A2(n762), .B1(n751), .B2(n777), .ZN(\U8/Z_19 )
         );
  INV_X4 U203 ( .A(n104), .ZN(\U8/Z_18 ) );
  INV_X4 U205 ( .A(n105), .ZN(\U8/Z_17 ) );
  OAI22_X2 U207 ( .A1(n724), .A2(n763), .B1(n751), .B2(n778), .ZN(\U8/Z_16 )
         );
  OAI22_X2 U210 ( .A1(n724), .A2(n764), .B1(n751), .B2(n779), .ZN(\U8/Z_15 )
         );
  OAI22_X2 U213 ( .A1(n724), .A2(n765), .B1(n751), .B2(n780), .ZN(\U8/Z_14 )
         );
  OAI22_X2 U216 ( .A1(n724), .A2(n766), .B1(n751), .B2(n781), .ZN(\U8/Z_13 )
         );
  INV_X4 U219 ( .A(n108), .ZN(\U8/Z_12 ) );
  INV_X4 U221 ( .A(n109), .ZN(\U8/Z_11 ) );
  OAI22_X2 U223 ( .A1(n724), .A2(n767), .B1(n751), .B2(n782), .ZN(\U8/Z_10 )
         );
  OAI22_X2 U226 ( .A1(n724), .A2(n773), .B1(n751), .B2(n788), .ZN(\U8/Z_1 ) );
  OAI22_X2 U229 ( .A1(n724), .A2(n774), .B1(n751), .B2(n789), .ZN(\U8/Z_0 ) );
  INV_X4 U232 ( .A(n111), .ZN(\U7/Z_9 ) );
  INV_X4 U234 ( .A(n112), .ZN(\U7/Z_8 ) );
  INV_X4 U236 ( .A(n113), .ZN(\U7/Z_7 ) );
  INV_X4 U238 ( .A(n114), .ZN(\U7/Z_6 ) );
  INV_X4 U240 ( .A(n115), .ZN(\U7/Z_5 ) );
  INV_X4 U242 ( .A(n116), .ZN(\U7/Z_4 ) );
  INV_X4 U244 ( .A(n117), .ZN(\U7/Z_3 ) );
  INV_X4 U246 ( .A(n118), .ZN(\U7/Z_23 ) );
  INV_X4 U248 ( .A(n119), .ZN(\U7/Z_22 ) );
  INV_X4 U250 ( .A(n120), .ZN(\U7/Z_21 ) );
  INV_X4 U252 ( .A(n121), .ZN(\U7/Z_20 ) );
  INV_X4 U254 ( .A(n122), .ZN(\U7/Z_2 ) );
  INV_X4 U256 ( .A(n123), .ZN(\U7/Z_19 ) );
  INV_X4 U258 ( .A(n124), .ZN(\U7/Z_18 ) );
  INV_X4 U260 ( .A(n125), .ZN(\U7/Z_17 ) );
  INV_X4 U262 ( .A(n126), .ZN(\U7/Z_16 ) );
  INV_X4 U264 ( .A(n127), .ZN(\U7/Z_15 ) );
  INV_X4 U266 ( .A(n128), .ZN(\U7/Z_14 ) );
  INV_X4 U268 ( .A(n129), .ZN(\U7/Z_13 ) );
  INV_X4 U270 ( .A(n130), .ZN(\U7/Z_12 ) );
  INV_X4 U272 ( .A(n131), .ZN(\U7/Z_11 ) );
  INV_X4 U274 ( .A(n132), .ZN(\U7/Z_10 ) );
  INV_X4 U276 ( .A(n133), .ZN(\U7/Z_1 ) );
  INV_X4 U278 ( .A(n134), .ZN(\U7/Z_0 ) );
  XOR2_X2 U282 ( .A(n384), .B(n385), .Z(n135) );
  NAND2_X2 U283 ( .A1(n136), .A2(n137), .ZN(\U4/Z_9 ) );
  NAND2_X2 U286 ( .A1(n142), .A2(n143), .ZN(\U4/Z_8 ) );
  NAND2_X2 U289 ( .A1(n144), .A2(n145), .ZN(\U4/Z_7 ) );
  NAND2_X2 U292 ( .A1(n146), .A2(n147), .ZN(\U4/Z_6 ) );
  NAND2_X2 U295 ( .A1(n148), .A2(n149), .ZN(\U4/Z_5 ) );
  NAND2_X2 U298 ( .A1(n150), .A2(n151), .ZN(\U4/Z_4 ) );
  NAND2_X2 U301 ( .A1(n152), .A2(n153), .ZN(\U4/Z_3 ) );
  NAND2_X2 U304 ( .A1(n154), .A2(n155), .ZN(\U4/Z_23 ) );
  NAND2_X2 U307 ( .A1(n156), .A2(n157), .ZN(\U4/Z_22 ) );
  NAND2_X2 U310 ( .A1(n158), .A2(n159), .ZN(\U4/Z_21 ) );
  NAND2_X2 U313 ( .A1(n160), .A2(n161), .ZN(\U4/Z_20 ) );
  NAND2_X2 U316 ( .A1(n162), .A2(n163), .ZN(\U4/Z_2 ) );
  NAND2_X2 U319 ( .A1(n164), .A2(n165), .ZN(\U4/Z_19 ) );
  NAND2_X2 U322 ( .A1(n166), .A2(n167), .ZN(\U4/Z_18 ) );
  NAND2_X2 U325 ( .A1(n168), .A2(n169), .ZN(\U4/Z_17 ) );
  NAND2_X2 U328 ( .A1(n170), .A2(n171), .ZN(\U4/Z_16 ) );
  NAND2_X2 U331 ( .A1(n172), .A2(n173), .ZN(\U4/Z_15 ) );
  NAND2_X2 U334 ( .A1(n174), .A2(n175), .ZN(\U4/Z_14 ) );
  NAND2_X2 U337 ( .A1(n176), .A2(n177), .ZN(\U4/Z_13 ) );
  NAND2_X2 U340 ( .A1(n178), .A2(n179), .ZN(\U4/Z_12 ) );
  NAND2_X2 U343 ( .A1(n180), .A2(n181), .ZN(\U4/Z_11 ) );
  NAND2_X2 U346 ( .A1(n182), .A2(n183), .ZN(\U4/Z_10 ) );
  NAND2_X2 U349 ( .A1(n184), .A2(n185), .ZN(\U4/Z_1 ) );
  NAND2_X2 U352 ( .A1(n186), .A2(n187), .ZN(\U4/Z_0 ) );
  AND4_X2 U355 ( .A1(n383), .A2(n32), .A3(\add_41/A[0] ), .A4(\add_41/A[1] ), 
        .ZN(n139) );
  AND4_X2 U358 ( .A1(n383), .A2(n32), .A3(n386), .A4(\add_41/A[1] ), .ZN(n141)
         );
  NOR2_X2 U360 ( .A1(n758), .A2(n384), .ZN(n32) );
  NOR3_X2 U362 ( .A1(\add_41/A[2] ), .A2(n383), .A3(n758), .ZN(n35) );
  DFF_X2 \Count_reg[4]  ( .D(n387), .CK(clock), .Q(n758), .QN(n382) );
  INV_X4 U27 ( .A(1'b0), .ZN(DiagonalYDone) );
  AND4_X4 U53 ( .A1(n32), .A2(n385), .A3(n386), .A4(\add_41/A[3] ), .ZN(n28)
         );
  NOR3_X2 U54 ( .A1(n720), .A2(reset), .A3(EnableChange), .ZN(n726) );
  AND4_X4 U79 ( .A1(n383), .A2(n386), .A3(n382), .A4(n135), .ZN(n724) );
  AND3_X4 U80 ( .A1(n386), .A2(n35), .A3(n385), .ZN(n721) );
  NOR3_X2 U82 ( .A1(n721), .A2(n141), .A3(n139), .ZN(n722) );
  INV_X4 U84 ( .A(n724), .ZN(n751) );
  INV_X4 U86 ( .A(n723), .ZN(n753) );
  INV_X4 U88 ( .A(n755), .ZN(n754) );
  AND3_X2 U90 ( .A1(\add_41/A[0] ), .A2(\add_41/A[1] ), .A3(n35), .ZN(n723) );
  INV_X4 U92 ( .A(n725), .ZN(n752) );
  INV_X4 U94 ( .A(n28), .ZN(n755) );
  INV_X4 U96 ( .A(n1), .ZN(n756) );
  AOI22_X2 U98 ( .A1(\U4/DATA1_0 ), .A2(n721), .B1(\U6/DATA1_0 ), .B2(n141), 
        .ZN(n186) );
  AOI22_X2 U100 ( .A1(\U6/DATA2_0 ), .A2(n722), .B1(\U5/DATA1_0 ), .B2(n139), 
        .ZN(n187) );
  AOI22_X2 U102 ( .A1(\U4/DATA1_1 ), .A2(n721), .B1(\U6/DATA1_1 ), .B2(n141), 
        .ZN(n184) );
  AOI22_X2 U104 ( .A1(\U6/DATA2_1 ), .A2(n722), .B1(\U5/DATA1_1 ), .B2(n139), 
        .ZN(n185) );
  AOI22_X2 U106 ( .A1(\U4/DATA1_2 ), .A2(n721), .B1(\U6/DATA1_2 ), .B2(n141), 
        .ZN(n162) );
  AOI22_X2 U108 ( .A1(\U6/DATA2_2 ), .A2(n722), .B1(\U5/DATA1_2 ), .B2(n139), 
        .ZN(n163) );
  AOI22_X2 U110 ( .A1(\U4/DATA1_3 ), .A2(n721), .B1(\U6/DATA1_3 ), .B2(n141), 
        .ZN(n152) );
  AOI22_X2 U112 ( .A1(\U6/DATA2_3 ), .A2(n722), .B1(\U5/DATA1_3 ), .B2(n139), 
        .ZN(n153) );
  AOI22_X2 U114 ( .A1(\U4/DATA1_4 ), .A2(n721), .B1(\U6/DATA1_4 ), .B2(n141), 
        .ZN(n150) );
  AOI22_X2 U116 ( .A1(\U6/DATA2_4 ), .A2(n722), .B1(\U5/DATA1_4 ), .B2(n139), 
        .ZN(n151) );
  AOI22_X2 U118 ( .A1(\U4/DATA1_5 ), .A2(n721), .B1(\U6/DATA1_5 ), .B2(n141), 
        .ZN(n148) );
  AOI22_X2 U120 ( .A1(\U6/DATA2_5 ), .A2(n722), .B1(\U5/DATA1_5 ), .B2(n139), 
        .ZN(n149) );
  AOI22_X2 U122 ( .A1(\U4/DATA1_6 ), .A2(n721), .B1(\U6/DATA1_6 ), .B2(n141), 
        .ZN(n146) );
  AOI22_X2 U124 ( .A1(\U6/DATA2_6 ), .A2(n722), .B1(\U5/DATA1_6 ), .B2(n139), 
        .ZN(n147) );
  AOI22_X2 U126 ( .A1(\U4/DATA1_7 ), .A2(n721), .B1(\U6/DATA1_7 ), .B2(n141), 
        .ZN(n144) );
  AOI22_X2 U128 ( .A1(\U6/DATA2_7 ), .A2(n722), .B1(\U5/DATA1_7 ), .B2(n139), 
        .ZN(n145) );
  AOI22_X2 U129 ( .A1(\U4/DATA1_8 ), .A2(n721), .B1(\U6/DATA1_8 ), .B2(n141), 
        .ZN(n142) );
  AOI22_X2 U130 ( .A1(\U6/DATA2_8 ), .A2(n722), .B1(\U5/DATA1_8 ), .B2(n139), 
        .ZN(n143) );
  AOI22_X2 U131 ( .A1(\U4/DATA1_9 ), .A2(n721), .B1(\U6/DATA1_9 ), .B2(n141), 
        .ZN(n136) );
  AOI22_X2 U132 ( .A1(\U6/DATA2_9 ), .A2(n722), .B1(\U5/DATA1_9 ), .B2(n139), 
        .ZN(n137) );
  AOI22_X2 U133 ( .A1(\U4/DATA1_10 ), .A2(n721), .B1(\U6/DATA1_10 ), .B2(n141), 
        .ZN(n182) );
  AOI22_X2 U137 ( .A1(\U6/DATA2_10 ), .A2(n722), .B1(\U5/DATA1_10 ), .B2(n139), 
        .ZN(n183) );
  AOI22_X2 U139 ( .A1(\U4/DATA1_11 ), .A2(n721), .B1(\U6/DATA1_11 ), .B2(n141), 
        .ZN(n180) );
  AOI22_X2 U141 ( .A1(\U6/DATA2_11 ), .A2(n722), .B1(\U5/DATA1_11 ), .B2(n139), 
        .ZN(n181) );
  AOI22_X2 U143 ( .A1(\U4/DATA1_12 ), .A2(n721), .B1(\U6/DATA1_12 ), .B2(n141), 
        .ZN(n178) );
  AOI22_X2 U145 ( .A1(\U6/DATA2_12 ), .A2(n722), .B1(\U5/DATA1_12 ), .B2(n139), 
        .ZN(n179) );
  AOI22_X2 U146 ( .A1(\U4/DATA1_13 ), .A2(n721), .B1(\U6/DATA1_13 ), .B2(n141), 
        .ZN(n176) );
  AOI22_X2 U148 ( .A1(\U6/DATA2_13 ), .A2(n722), .B1(\U5/DATA1_13 ), .B2(n139), 
        .ZN(n177) );
  AOI22_X2 U162 ( .A1(\U4/DATA1_14 ), .A2(n721), .B1(\U6/DATA1_14 ), .B2(n141), 
        .ZN(n174) );
  AOI22_X2 U170 ( .A1(\U6/DATA2_14 ), .A2(n722), .B1(\U5/DATA1_14 ), .B2(n139), 
        .ZN(n175) );
  AOI22_X2 U172 ( .A1(\U4/DATA1_15 ), .A2(n721), .B1(\U6/DATA1_15 ), .B2(n141), 
        .ZN(n172) );
  AOI22_X2 U174 ( .A1(\U6/DATA2_15 ), .A2(n722), .B1(\U5/DATA1_15 ), .B2(n139), 
        .ZN(n173) );
  AOI22_X2 U176 ( .A1(\U4/DATA1_16 ), .A2(n721), .B1(\U6/DATA1_16 ), .B2(n141), 
        .ZN(n170) );
  AOI22_X2 U177 ( .A1(\U6/DATA2_16 ), .A2(n722), .B1(\U5/DATA1_16 ), .B2(n139), 
        .ZN(n171) );
  AOI22_X2 U179 ( .A1(\U4/DATA1_17 ), .A2(n721), .B1(\U6/DATA1_17 ), .B2(n141), 
        .ZN(n168) );
  AOI22_X2 U180 ( .A1(\U6/DATA2_17 ), .A2(n722), .B1(\U5/DATA1_17 ), .B2(n139), 
        .ZN(n169) );
  AOI22_X2 U182 ( .A1(\U4/DATA1_18 ), .A2(n721), .B1(\U6/DATA1_18 ), .B2(n141), 
        .ZN(n166) );
  AOI22_X2 U183 ( .A1(\U6/DATA2_18 ), .A2(n722), .B1(\U5/DATA1_18 ), .B2(n139), 
        .ZN(n167) );
  AOI22_X2 U185 ( .A1(\U4/DATA1_19 ), .A2(n721), .B1(\U6/DATA1_19 ), .B2(n141), 
        .ZN(n164) );
  AOI22_X2 U186 ( .A1(\U6/DATA2_19 ), .A2(n722), .B1(\U5/DATA1_19 ), .B2(n139), 
        .ZN(n165) );
  AOI22_X2 U188 ( .A1(\U4/DATA1_20 ), .A2(n721), .B1(\U6/DATA1_20 ), .B2(n141), 
        .ZN(n160) );
  AOI22_X2 U190 ( .A1(\U6/DATA2_20 ), .A2(n722), .B1(\U5/DATA1_20 ), .B2(n139), 
        .ZN(n161) );
  AOI22_X2 U192 ( .A1(\U4/DATA1_21 ), .A2(n721), .B1(\U6/DATA1_21 ), .B2(n141), 
        .ZN(n158) );
  AOI22_X2 U193 ( .A1(\U6/DATA2_21 ), .A2(n722), .B1(\U5/DATA1_21 ), .B2(n139), 
        .ZN(n159) );
  AOI22_X2 U195 ( .A1(\U4/DATA1_22 ), .A2(n721), .B1(\U6/DATA1_22 ), .B2(n141), 
        .ZN(n156) );
  AOI22_X2 U196 ( .A1(\U6/DATA2_22 ), .A2(n722), .B1(\U5/DATA1_22 ), .B2(n139), 
        .ZN(n157) );
  AOI22_X2 U198 ( .A1(\U4/DATA1_23 ), .A2(n721), .B1(\U6/DATA1_23 ), .B2(n141), 
        .ZN(n154) );
  AOI22_X2 U199 ( .A1(\U6/DATA2_23 ), .A2(n722), .B1(\U5/DATA1_23 ), .B2(n139), 
        .ZN(n155) );
  OAI21_X2 U201 ( .B1(n383), .B2(n47), .A(n48), .ZN(n388) );
  OAI21_X2 U202 ( .B1(n384), .B2(n47), .A(n49), .ZN(n389) );
  OAI21_X2 U204 ( .B1(n385), .B2(n47), .A(n50), .ZN(n390) );
  OAI21_X2 U206 ( .B1(n44), .B2(n759), .A(n758), .ZN(n41) );
  AOI22_X2 U208 ( .A1(\add_41/A[0] ), .A2(n759), .B1(n386), .B2(n43), .ZN(n51)
         );
  AOI22_X2 U209 ( .A1(\U11/DATA1_0 ), .A2(n724), .B1(\U11/DATA2_0 ), .B2(n751), 
        .ZN(n134) );
  AOI22_X2 U211 ( .A1(\U11/DATA1_1 ), .A2(n724), .B1(\U11/DATA2_1 ), .B2(n751), 
        .ZN(n133) );
  AOI22_X2 U212 ( .A1(\U11/DATA1_10 ), .A2(n724), .B1(\U11/DATA2_10 ), .B2(
        n751), .ZN(n132) );
  AOI22_X2 U214 ( .A1(\U11/DATA1_11 ), .A2(n724), .B1(\U11/DATA2_11 ), .B2(
        n751), .ZN(n131) );
  AOI22_X2 U215 ( .A1(\U11/DATA1_12 ), .A2(n724), .B1(\U11/DATA2_12 ), .B2(
        n751), .ZN(n130) );
  AOI22_X2 U217 ( .A1(\U11/DATA1_13 ), .A2(n724), .B1(\U11/DATA2_13 ), .B2(
        n751), .ZN(n129) );
  AOI22_X2 U218 ( .A1(\U11/DATA1_14 ), .A2(n724), .B1(\U11/DATA2_14 ), .B2(
        n751), .ZN(n128) );
  AOI22_X2 U220 ( .A1(\U11/DATA1_15 ), .A2(n724), .B1(\U11/DATA2_15 ), .B2(
        n751), .ZN(n127) );
  AOI22_X2 U222 ( .A1(\U11/DATA1_17 ), .A2(n724), .B1(\U11/DATA2_17 ), .B2(
        n751), .ZN(n125) );
  AOI22_X2 U224 ( .A1(\U11/DATA1_18 ), .A2(n724), .B1(\U11/DATA2_18 ), .B2(
        n751), .ZN(n124) );
  AOI22_X2 U225 ( .A1(\U11/DATA1_19 ), .A2(n724), .B1(\U11/DATA2_19 ), .B2(
        n751), .ZN(n123) );
  AOI22_X2 U227 ( .A1(\U11/DATA1_20 ), .A2(n724), .B1(\U11/DATA2_20 ), .B2(
        n751), .ZN(n121) );
  AOI22_X2 U228 ( .A1(n751), .A2(\U12/DATA2_7 ), .B1(n724), .B2(\U12/DATA1_7 ), 
        .ZN(n97) );
  AOI22_X2 U230 ( .A1(n751), .A2(\U12/DATA2_8 ), .B1(n724), .B2(\U12/DATA1_8 ), 
        .ZN(n96) );
  AOI22_X2 U231 ( .A1(n751), .A2(\U12/DATA2_9 ), .B1(n724), .B2(\U12/DATA1_9 ), 
        .ZN(n93) );
  AOI22_X2 U233 ( .A1(n751), .A2(\U12/DATA2_11 ), .B1(n724), .B2(
        \U12/DATA1_11 ), .ZN(n109) );
  AOI22_X2 U235 ( .A1(n751), .A2(\U12/DATA2_22 ), .B1(n724), .B2(
        \U12/DATA1_22 ), .ZN(n101) );
  AOI22_X2 U237 ( .A1(\U11/DATA1_2 ), .A2(n724), .B1(\U11/DATA2_2 ), .B2(n751), 
        .ZN(n122) );
  AOI22_X2 U239 ( .A1(\U11/DATA1_3 ), .A2(n724), .B1(\U11/DATA2_3 ), .B2(n751), 
        .ZN(n117) );
  AOI22_X2 U241 ( .A1(\U11/DATA1_4 ), .A2(n724), .B1(\U11/DATA2_4 ), .B2(n751), 
        .ZN(n116) );
  AOI22_X2 U243 ( .A1(\U11/DATA1_5 ), .A2(n724), .B1(\U11/DATA2_5 ), .B2(n751), 
        .ZN(n115) );
  AOI22_X2 U245 ( .A1(\U11/DATA1_6 ), .A2(n724), .B1(\U11/DATA2_6 ), .B2(n751), 
        .ZN(n114) );
  AOI22_X2 U247 ( .A1(\U11/DATA1_7 ), .A2(n724), .B1(\U11/DATA2_7 ), .B2(n751), 
        .ZN(n113) );
  AOI22_X2 U249 ( .A1(\U11/DATA1_8 ), .A2(n724), .B1(\U11/DATA2_8 ), .B2(n751), 
        .ZN(n112) );
  AOI22_X2 U251 ( .A1(\U11/DATA1_9 ), .A2(n724), .B1(\U11/DATA2_9 ), .B2(n751), 
        .ZN(n111) );
  AOI22_X2 U253 ( .A1(\U11/DATA1_16 ), .A2(n724), .B1(\U11/DATA2_16 ), .B2(
        n751), .ZN(n126) );
  AOI22_X2 U255 ( .A1(\U11/DATA1_21 ), .A2(n724), .B1(\U11/DATA2_21 ), .B2(
        n751), .ZN(n120) );
  AOI22_X2 U257 ( .A1(\U11/DATA1_22 ), .A2(n724), .B1(\U11/DATA2_22 ), .B2(
        n751), .ZN(n119) );
  AOI22_X2 U259 ( .A1(\U11/DATA1_23 ), .A2(n724), .B1(\U11/DATA2_23 ), .B2(
        n751), .ZN(n118) );
  AOI22_X2 U261 ( .A1(n751), .A2(\U12/DATA2_12 ), .B1(n724), .B2(
        \U12/DATA1_12 ), .ZN(n108) );
  AOI22_X2 U263 ( .A1(n751), .A2(\U12/DATA2_17 ), .B1(n724), .B2(
        \U12/DATA1_17 ), .ZN(n105) );
  AOI22_X2 U265 ( .A1(n751), .A2(\U12/DATA2_18 ), .B1(n724), .B2(
        \U12/DATA1_18 ), .ZN(n104) );
  AOI22_X2 U267 ( .A1(n751), .A2(\U12/DATA2_23 ), .B1(n724), .B2(
        \U12/DATA1_23 ), .ZN(n100) );
  AND3_X2 U269 ( .A1(n35), .A2(\add_41/A[0] ), .A3(n385), .ZN(n725) );
  OR2_X1 U271 ( .A1(n756), .A2(n726), .ZN(n381) );
  BUF_X4 U273 ( .A(SubOutput[0]), .Z(AddInput2[0]) );
  BUF_X4 U275 ( .A(SubOutput[1]), .Z(AddInput2[1]) );
  BUF_X4 U277 ( .A(SubOutput[2]), .Z(AddInput2[2]) );
  BUF_X4 U279 ( .A(SubOutput[3]), .Z(AddInput2[3]) );
  BUF_X4 U280 ( .A(SubOutput[4]), .Z(AddInput2[4]) );
  BUF_X4 U281 ( .A(SubOutput[5]), .Z(AddInput2[5]) );
  BUF_X4 U284 ( .A(SubOutput[6]), .Z(AddInput2[6]) );
  BUF_X4 U285 ( .A(SubOutput[7]), .Z(AddInput2[7]) );
  BUF_X4 U287 ( .A(SubOutput[8]), .Z(AddInput2[8]) );
  BUF_X4 U288 ( .A(SubOutput[9]), .Z(AddInput2[9]) );
  BUF_X4 U290 ( .A(SubOutput[10]), .Z(AddInput2[10]) );
  BUF_X4 U291 ( .A(SubOutput[11]), .Z(AddInput2[11]) );
  BUF_X4 U293 ( .A(SubOutput[12]), .Z(AddInput2[12]) );
  BUF_X4 U294 ( .A(SubOutput[13]), .Z(AddInput2[13]) );
  BUF_X4 U296 ( .A(SubOutput[14]), .Z(AddInput2[14]) );
  BUF_X4 U297 ( .A(SubOutput[15]), .Z(AddInput2[15]) );
  BUF_X4 U299 ( .A(SubOutput[16]), .Z(AddInput2[16]) );
  BUF_X4 U300 ( .A(SubOutput[17]), .Z(AddInput2[17]) );
  BUF_X4 U302 ( .A(SubOutput[18]), .Z(AddInput2[18]) );
  BUF_X4 U303 ( .A(SubOutput[19]), .Z(AddInput2[19]) );
  BUF_X4 U305 ( .A(SubOutput[20]), .Z(AddInput2[20]) );
  BUF_X4 U306 ( .A(SubOutput[21]), .Z(AddInput2[21]) );
  BUF_X4 U308 ( .A(SubOutput[22]), .Z(AddInput2[22]) );
  BUF_X4 U309 ( .A(SubOutput[23]), .Z(AddInput2[23]) );
  INV_X4 U311 ( .A(n51), .ZN(n757) );
  INV_X4 U312 ( .A(n47), .ZN(n759) );
  INV_X4 U314 ( .A(\U12/DATA2_21 ), .ZN(n760) );
  INV_X4 U315 ( .A(\U12/DATA2_20 ), .ZN(n761) );
  INV_X4 U317 ( .A(\U12/DATA2_19 ), .ZN(n762) );
  INV_X4 U318 ( .A(\U12/DATA2_16 ), .ZN(n763) );
  INV_X4 U320 ( .A(\U12/DATA2_15 ), .ZN(n764) );
  INV_X4 U321 ( .A(\U12/DATA2_14 ), .ZN(n765) );
  INV_X4 U323 ( .A(\U12/DATA2_13 ), .ZN(n766) );
  INV_X4 U324 ( .A(\U12/DATA2_10 ), .ZN(n767) );
  INV_X4 U326 ( .A(\U12/DATA2_6 ), .ZN(n768) );
  INV_X4 U327 ( .A(\U12/DATA2_5 ), .ZN(n769) );
  INV_X4 U329 ( .A(\U12/DATA2_4 ), .ZN(n770) );
  INV_X4 U330 ( .A(\U12/DATA2_3 ), .ZN(n771) );
  INV_X4 U332 ( .A(\U12/DATA2_2 ), .ZN(n772) );
  INV_X4 U333 ( .A(\U12/DATA2_1 ), .ZN(n773) );
  INV_X4 U335 ( .A(\U12/DATA2_0 ), .ZN(n774) );
  INV_X4 U336 ( .A(\U12/DATA1_21 ), .ZN(n775) );
  INV_X4 U338 ( .A(\U12/DATA1_20 ), .ZN(n776) );
  INV_X4 U339 ( .A(\U12/DATA1_19 ), .ZN(n777) );
  INV_X4 U341 ( .A(\U12/DATA1_16 ), .ZN(n778) );
  INV_X4 U342 ( .A(\U12/DATA1_15 ), .ZN(n779) );
  INV_X4 U344 ( .A(\U12/DATA1_14 ), .ZN(n780) );
  INV_X4 U345 ( .A(\U12/DATA1_13 ), .ZN(n781) );
  INV_X4 U347 ( .A(\U12/DATA1_10 ), .ZN(n782) );
  INV_X4 U348 ( .A(\U12/DATA1_6 ), .ZN(n783) );
  INV_X4 U350 ( .A(\U12/DATA1_5 ), .ZN(n784) );
  INV_X4 U351 ( .A(\U12/DATA1_4 ), .ZN(n785) );
  INV_X4 U353 ( .A(\U12/DATA1_3 ), .ZN(n786) );
  INV_X4 U354 ( .A(\U12/DATA1_2 ), .ZN(n787) );
  INV_X4 U356 ( .A(\U12/DATA1_1 ), .ZN(n788) );
  INV_X4 U357 ( .A(\U12/DATA1_0 ), .ZN(n789) );
  INV_X4 U359 ( .A(EnableChange), .ZN(n790) );
  INV_X4 U361 ( .A(AddOutput[23]), .ZN(n791) );
  INV_X4 U363 ( .A(AddOutput[22]), .ZN(n792) );
  INV_X4 U364 ( .A(AddOutput[21]), .ZN(n793) );
  INV_X4 U366 ( .A(AddOutput[20]), .ZN(n794) );
  INV_X4 U367 ( .A(AddOutput[19]), .ZN(n795) );
  INV_X4 U368 ( .A(AddOutput[18]), .ZN(n796) );
  INV_X4 U369 ( .A(AddOutput[17]), .ZN(n797) );
  INV_X4 U370 ( .A(AddOutput[16]), .ZN(n798) );
  INV_X4 U371 ( .A(AddOutput[15]), .ZN(n799) );
  INV_X4 U372 ( .A(AddOutput[14]), .ZN(n800) );
  INV_X4 U373 ( .A(AddOutput[13]), .ZN(n801) );
  INV_X4 U374 ( .A(AddOutput[12]), .ZN(n802) );
  INV_X4 U375 ( .A(AddOutput[11]), .ZN(n803) );
  INV_X4 U376 ( .A(AddOutput[10]), .ZN(n804) );
  INV_X4 U377 ( .A(AddOutput[9]), .ZN(n805) );
  INV_X4 U378 ( .A(AddOutput[8]), .ZN(n806) );
  INV_X4 U379 ( .A(AddOutput[7]), .ZN(n807) );
  INV_X4 U380 ( .A(AddOutput[6]), .ZN(n808) );
  INV_X4 U381 ( .A(AddOutput[5]), .ZN(n809) );
  INV_X4 U382 ( .A(AddOutput[4]), .ZN(n810) );
  INV_X4 U383 ( .A(AddOutput[3]), .ZN(n811) );
  INV_X4 U384 ( .A(AddOutput[2]), .ZN(n812) );
  INV_X4 U385 ( .A(AddOutput[1]), .ZN(n813) );
  INV_X4 U386 ( .A(AddOutput[0]), .ZN(n814) );
endmodule


module pad_3 ( Element, PosElement, Y_ramRow, PaddedRow, RowReady );
  input [47:0] Element;
  input [12:0] PosElement;
  input [255:0] Y_ramRow;
  output [255:0] PaddedRow;
  output RowReady;
  wire   \U7/DATA1_0 , \U7/DATA1_1 , \U7/DATA1_2 , \U7/DATA1_3 , \U7/DATA1_4 ,
         \U7/DATA1_5 , \U7/DATA1_6 , \U7/DATA1_7 , \U7/DATA1_8 , \U7/DATA1_9 ,
         \U7/DATA1_10 , \U7/DATA1_11 , \U7/DATA1_12 , \U7/DATA1_13 ,
         \U7/DATA1_14 , \U7/DATA1_15 , \U7/DATA1_16 , \U7/DATA1_17 ,
         \U7/DATA1_18 , \U7/DATA1_19 , \U7/DATA1_20 , \U7/DATA1_21 ,
         \U7/DATA1_22 , \U7/DATA1_23 , \U7/DATA1_24 , \U7/DATA1_25 ,
         \U7/DATA1_26 , \U7/DATA1_27 , \U7/DATA1_28 , \U7/DATA1_29 ,
         \U7/DATA1_30 , \U7/DATA1_31 , \U7/DATA1_32 , \U7/DATA1_33 ,
         \U7/DATA1_34 , \U7/DATA1_35 , \U7/DATA1_36 , \U7/DATA1_37 ,
         \U7/DATA1_38 , \U7/DATA1_39 , \U7/DATA1_40 , \U7/DATA1_41 ,
         \U7/DATA1_42 , \U7/DATA1_43 , \U7/DATA1_44 , \U7/DATA1_45 ,
         \U7/DATA1_46 , \U7/DATA1_47 , \U7/DATA1_64 , \U7/DATA1_65 ,
         \U7/DATA1_66 , \U7/DATA1_67 , \U7/DATA1_68 , \U7/DATA1_69 ,
         \U7/DATA1_70 , \U7/DATA1_71 , \U7/DATA1_72 , \U7/DATA1_73 ,
         \U7/DATA1_74 , \U7/DATA1_75 , \U7/DATA1_76 , \U7/DATA1_77 ,
         \U7/DATA1_78 , \U7/DATA1_79 , \U7/DATA1_80 , \U7/DATA1_81 ,
         \U7/DATA1_82 , \U7/DATA1_83 , \U7/DATA1_84 , \U7/DATA1_85 ,
         \U7/DATA1_86 , \U7/DATA1_87 , \U7/DATA1_88 , \U7/DATA1_89 ,
         \U7/DATA1_90 , \U7/DATA1_91 , \U7/DATA1_92 , \U7/DATA1_93 ,
         \U7/DATA1_94 , \U7/DATA1_95 , \U7/DATA1_96 , \U7/DATA1_97 ,
         \U7/DATA1_98 , \U7/DATA1_99 , \U7/DATA1_100 , \U7/DATA1_101 ,
         \U7/DATA1_102 , \U7/DATA1_103 , \U7/DATA1_104 , \U7/DATA1_105 ,
         \U7/DATA1_106 , \U7/DATA1_107 , \U7/DATA1_108 , \U7/DATA1_109 ,
         \U7/DATA1_110 , \U7/DATA1_111 , \U7/DATA1_128 , \U7/DATA1_129 ,
         \U7/DATA1_130 , \U7/DATA1_131 , \U7/DATA1_132 , \U7/DATA1_133 ,
         \U7/DATA1_134 , \U7/DATA1_135 , \U7/DATA1_136 , \U7/DATA1_137 ,
         \U7/DATA1_138 , \U7/DATA1_139 , \U7/DATA1_140 , \U7/DATA1_141 ,
         \U7/DATA1_142 , \U7/DATA1_143 , \U7/DATA1_144 , \U7/DATA1_145 ,
         \U7/DATA1_146 , \U7/DATA1_147 , \U7/DATA1_148 , \U7/DATA1_149 ,
         \U7/DATA1_150 , \U7/DATA1_151 , \U7/DATA1_152 , \U7/DATA1_153 ,
         \U7/DATA1_154 , \U7/DATA1_155 , \U7/DATA1_156 , \U7/DATA1_157 ,
         \U7/DATA1_158 , \U7/DATA1_159 , \U7/DATA1_160 , \U7/DATA1_161 ,
         \U7/DATA1_162 , \U7/DATA1_163 , \U7/DATA1_164 , \U7/DATA1_165 ,
         \U7/DATA1_166 , \U7/DATA1_167 , \U7/DATA1_168 , \U7/DATA1_169 ,
         \U7/DATA1_170 , \U7/DATA1_171 , \U7/DATA1_172 , \U7/DATA1_173 ,
         \U7/DATA1_174 , \U7/DATA1_175 , \U7/DATA1_192 , \U7/DATA1_193 ,
         \U7/DATA1_194 , \U7/DATA1_195 , \U7/DATA1_196 , \U7/DATA1_197 ,
         \U7/DATA1_198 , \U7/DATA1_199 , \U7/DATA1_200 , \U7/DATA1_201 ,
         \U7/DATA1_202 , \U7/DATA1_203 , \U7/DATA1_204 , \U7/DATA1_205 ,
         \U7/DATA1_206 , \U7/DATA1_207 , \U7/DATA1_208 , \U7/DATA1_209 ,
         \U7/DATA1_210 , \U7/DATA1_211 , \U7/DATA1_212 , \U7/DATA1_213 ,
         \U7/DATA1_214 , \U7/DATA1_215 , \U7/DATA1_216 , \U7/DATA1_217 ,
         \U7/DATA1_218 , \U7/DATA1_219 , \U7/DATA1_220 , \U7/DATA1_221 ,
         \U7/DATA1_222 , \U7/DATA1_223 , \U7/DATA1_224 , \U7/DATA1_225 ,
         \U7/DATA1_226 , \U7/DATA1_227 , \U7/DATA1_228 , \U7/DATA1_229 ,
         \U7/DATA1_230 , \U7/DATA1_231 , \U7/DATA1_232 , \U7/DATA1_233 ,
         \U7/DATA1_234 , \U7/DATA1_235 , \U7/DATA1_236 , \U7/DATA1_237 ,
         \U7/DATA1_238 , \U7/DATA1_239 , \U6/DATA1_192 , \U6/DATA1_193 ,
         \U6/DATA1_194 , \U6/DATA1_195 , \U6/DATA1_196 , \U6/DATA1_197 ,
         \U6/DATA1_198 , \U6/DATA1_199 , \U6/DATA1_200 , \U6/DATA1_201 ,
         \U6/DATA1_202 , \U6/DATA1_203 , \U6/DATA1_204 , \U6/DATA1_205 ,
         \U6/DATA1_206 , \U6/DATA1_207 , \U6/DATA1_208 , \U6/DATA1_209 ,
         \U6/DATA1_210 , \U6/DATA1_211 , \U6/DATA1_212 , \U6/DATA1_213 ,
         \U6/DATA1_214 , \U6/DATA1_215 , \U6/DATA1_216 , \U6/DATA1_217 ,
         \U6/DATA1_218 , \U6/DATA1_219 , \U6/DATA1_220 , \U6/DATA1_221 ,
         \U6/DATA1_222 , \U6/DATA1_223 , \U6/DATA1_224 , \U6/DATA1_225 ,
         \U6/DATA1_226 , \U6/DATA1_227 , \U6/DATA1_228 , \U6/DATA1_229 ,
         \U6/DATA1_230 , \U6/DATA1_231 , \U6/DATA1_232 , \U6/DATA1_233 ,
         \U6/DATA1_234 , \U6/DATA1_235 , \U6/DATA1_236 , \U6/DATA1_237 ,
         \U6/DATA1_238 , \U6/DATA1_239 , \U4/Z_0 , \U4/Z_1 , \U4/Z_2 ,
         \U4/Z_3 , \U4/Z_4 , \U4/Z_5 , \U4/Z_6 , \U4/Z_7 , \U4/Z_8 , \U4/Z_9 ,
         \U4/Z_10 , \U4/Z_11 , \U4/Z_12 , \U4/Z_13 , \U4/Z_14 , \U4/Z_15 ,
         \U4/Z_16 , \U4/Z_17 , \U4/Z_18 , \U4/Z_19 , \U4/Z_20 , \U4/Z_21 ,
         \U4/Z_22 , \U4/Z_23 , \U4/Z_24 , \U4/Z_25 , \U4/Z_26 , \U4/Z_27 ,
         \U4/Z_28 , \U4/Z_29 , \U4/Z_30 , \U4/Z_31 , \U4/Z_32 , \U4/Z_33 ,
         \U4/Z_34 , \U4/Z_35 , \U4/Z_36 , \U4/Z_37 , \U4/Z_38 , \U4/Z_39 ,
         \U4/Z_40 , \U4/Z_41 , \U4/Z_42 , \U4/Z_43 , \U4/Z_44 , \U4/Z_45 ,
         \U4/Z_46 , \U4/Z_47 , \U4/Z_48 , \U4/Z_49 , \U4/Z_50 , \U4/Z_51 ,
         \U4/Z_52 , \U4/Z_53 , \U4/Z_54 , \U4/Z_55 , \U4/Z_56 , \U4/Z_57 ,
         \U4/Z_58 , \U4/Z_59 , \U4/Z_60 , \U4/Z_61 , \U4/Z_62 , \U4/Z_63 ,
         \U4/Z_64 , \U4/Z_65 , \U4/Z_66 , \U4/Z_67 , \U4/Z_68 , \U4/Z_69 ,
         \U4/Z_70 , \U4/Z_71 , \U4/Z_72 , \U4/Z_73 , \U4/Z_74 , \U4/Z_75 ,
         \U4/Z_76 , \U4/Z_77 , \U4/Z_78 , \U4/Z_79 , \U4/Z_80 , \U4/Z_81 ,
         \U4/Z_82 , \U4/Z_83 , \U4/Z_84 , \U4/Z_85 , \U4/Z_86 , \U4/Z_87 ,
         \U4/Z_88 , \U4/Z_89 , \U4/Z_90 , \U4/Z_91 , \U4/Z_92 , \U4/Z_93 ,
         \U4/Z_94 , \U4/Z_95 , \U4/Z_96 , \U4/Z_97 , \U4/Z_98 , \U4/Z_99 ,
         \U4/Z_100 , \U4/Z_101 , \U4/Z_102 , \U4/Z_103 , \U4/Z_104 ,
         \U4/Z_105 , \U4/Z_106 , \U4/Z_107 , \U4/Z_108 , \U4/Z_109 ,
         \U4/Z_110 , \U4/Z_111 , \U4/Z_112 , \U4/Z_113 , \U4/Z_114 ,
         \U4/Z_115 , \U4/Z_116 , \U4/Z_117 , \U4/Z_118 , \U4/Z_119 ,
         \U4/Z_120 , \U4/Z_121 , \U4/Z_122 , \U4/Z_123 , \U4/Z_124 ,
         \U4/Z_125 , \U4/Z_126 , \U4/Z_127 , \U4/Z_128 , \U4/Z_129 ,
         \U4/Z_130 , \U4/Z_131 , \U4/Z_132 , \U4/Z_133 , \U4/Z_134 ,
         \U4/Z_135 , \U4/Z_136 , \U4/Z_137 , \U4/Z_138 , \U4/Z_139 ,
         \U4/Z_140 , \U4/Z_141 , \U4/Z_142 , \U4/Z_143 , \U4/Z_144 ,
         \U4/Z_145 , \U4/Z_146 , \U4/Z_147 , \U4/Z_148 , \U4/Z_149 ,
         \U4/Z_150 , \U4/Z_151 , \U4/Z_152 , \U4/Z_153 , \U4/Z_154 ,
         \U4/Z_155 , \U4/Z_156 , \U4/Z_157 , \U4/Z_158 , \U4/Z_159 ,
         \U4/Z_160 , \U4/Z_161 , \U4/Z_162 , \U4/Z_163 , \U4/Z_164 ,
         \U4/Z_165 , \U4/Z_166 , \U4/Z_167 , \U4/Z_168 , \U4/Z_169 ,
         \U4/Z_170 , \U4/Z_171 , \U4/Z_172 , \U4/Z_173 , \U4/Z_174 ,
         \U4/Z_175 , \U4/Z_176 , \U4/Z_177 , \U4/Z_178 , \U4/Z_179 ,
         \U4/Z_180 , \U4/Z_181 , \U4/Z_182 , \U4/Z_183 , \U4/Z_184 ,
         \U4/Z_185 , \U4/Z_186 , \U4/Z_187 , \U4/Z_188 , \U4/Z_189 ,
         \U4/Z_190 , \U4/Z_191 , \U4/Z_192 , \U4/Z_193 , \U4/Z_194 ,
         \U4/Z_195 , \U4/Z_196 , \U4/Z_197 , \U4/Z_198 , \U4/Z_199 ,
         \U4/Z_200 , \U4/Z_201 , \U4/Z_202 , \U4/Z_203 , \U4/Z_204 ,
         \U4/Z_205 , \U4/Z_206 , \U4/Z_207 , \U4/Z_208 , \U4/Z_209 ,
         \U4/Z_210 , \U4/Z_211 , \U4/Z_212 , \U4/Z_213 , \U4/Z_214 ,
         \U4/Z_215 , \U4/Z_216 , \U4/Z_217 , \U4/Z_218 , \U4/Z_219 ,
         \U4/Z_220 , \U4/Z_221 , \U4/Z_222 , \U4/Z_223 , \U4/Z_224 ,
         \U4/Z_225 , \U4/Z_226 , \U4/Z_227 , \U4/Z_228 , \U4/Z_229 ,
         \U4/Z_230 , \U4/Z_231 , \U4/Z_232 , \U4/Z_233 , \U4/Z_234 ,
         \U4/Z_235 , \U4/Z_236 , \U4/Z_237 , \U4/Z_238 , \U4/Z_239 ,
         \U4/Z_240 , \U4/Z_241 , \U4/Z_242 , \U4/Z_243 , \U4/Z_244 ,
         \U4/Z_245 , \U4/Z_246 , \U4/Z_247 , \U4/Z_248 , \U4/Z_249 ,
         \U4/Z_250 , \U4/Z_251 , \U4/Z_252 , \U4/Z_253 , \U4/Z_254 ,
         \U4/Z_255 , n50, n51, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n1363, n1364, n1365, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485;
  assign \U7/DATA1_0  = Y_ramRow[0];
  assign \U7/DATA1_1  = Y_ramRow[1];
  assign \U7/DATA1_2  = Y_ramRow[2];
  assign \U7/DATA1_3  = Y_ramRow[3];
  assign \U7/DATA1_4  = Y_ramRow[4];
  assign \U7/DATA1_5  = Y_ramRow[5];
  assign \U7/DATA1_6  = Y_ramRow[6];
  assign \U7/DATA1_7  = Y_ramRow[7];
  assign \U7/DATA1_8  = Y_ramRow[8];
  assign \U7/DATA1_9  = Y_ramRow[9];
  assign \U7/DATA1_10  = Y_ramRow[10];
  assign \U7/DATA1_11  = Y_ramRow[11];
  assign \U7/DATA1_12  = Y_ramRow[12];
  assign \U7/DATA1_13  = Y_ramRow[13];
  assign \U7/DATA1_14  = Y_ramRow[14];
  assign \U7/DATA1_15  = Y_ramRow[15];
  assign \U7/DATA1_16  = Y_ramRow[16];
  assign \U7/DATA1_17  = Y_ramRow[17];
  assign \U7/DATA1_18  = Y_ramRow[18];
  assign \U7/DATA1_19  = Y_ramRow[19];
  assign \U7/DATA1_20  = Y_ramRow[20];
  assign \U7/DATA1_21  = Y_ramRow[21];
  assign \U7/DATA1_22  = Y_ramRow[22];
  assign \U7/DATA1_23  = Y_ramRow[23];
  assign \U7/DATA1_24  = Y_ramRow[24];
  assign \U7/DATA1_25  = Y_ramRow[25];
  assign \U7/DATA1_26  = Y_ramRow[26];
  assign \U7/DATA1_27  = Y_ramRow[27];
  assign \U7/DATA1_28  = Y_ramRow[28];
  assign \U7/DATA1_29  = Y_ramRow[29];
  assign \U7/DATA1_30  = Y_ramRow[30];
  assign \U7/DATA1_31  = Y_ramRow[31];
  assign \U7/DATA1_32  = Y_ramRow[32];
  assign \U7/DATA1_33  = Y_ramRow[33];
  assign \U7/DATA1_34  = Y_ramRow[34];
  assign \U7/DATA1_35  = Y_ramRow[35];
  assign \U7/DATA1_36  = Y_ramRow[36];
  assign \U7/DATA1_37  = Y_ramRow[37];
  assign \U7/DATA1_38  = Y_ramRow[38];
  assign \U7/DATA1_39  = Y_ramRow[39];
  assign \U7/DATA1_40  = Y_ramRow[40];
  assign \U7/DATA1_41  = Y_ramRow[41];
  assign \U7/DATA1_42  = Y_ramRow[42];
  assign \U7/DATA1_43  = Y_ramRow[43];
  assign \U7/DATA1_44  = Y_ramRow[44];
  assign \U7/DATA1_45  = Y_ramRow[45];
  assign \U7/DATA1_46  = Y_ramRow[46];
  assign \U7/DATA1_47  = Y_ramRow[47];
  assign \U7/DATA1_64  = Y_ramRow[64];
  assign \U7/DATA1_65  = Y_ramRow[65];
  assign \U7/DATA1_66  = Y_ramRow[66];
  assign \U7/DATA1_67  = Y_ramRow[67];
  assign \U7/DATA1_68  = Y_ramRow[68];
  assign \U7/DATA1_69  = Y_ramRow[69];
  assign \U7/DATA1_70  = Y_ramRow[70];
  assign \U7/DATA1_71  = Y_ramRow[71];
  assign \U7/DATA1_72  = Y_ramRow[72];
  assign \U7/DATA1_73  = Y_ramRow[73];
  assign \U7/DATA1_74  = Y_ramRow[74];
  assign \U7/DATA1_75  = Y_ramRow[75];
  assign \U7/DATA1_76  = Y_ramRow[76];
  assign \U7/DATA1_77  = Y_ramRow[77];
  assign \U7/DATA1_78  = Y_ramRow[78];
  assign \U7/DATA1_79  = Y_ramRow[79];
  assign \U7/DATA1_80  = Y_ramRow[80];
  assign \U7/DATA1_81  = Y_ramRow[81];
  assign \U7/DATA1_82  = Y_ramRow[82];
  assign \U7/DATA1_83  = Y_ramRow[83];
  assign \U7/DATA1_84  = Y_ramRow[84];
  assign \U7/DATA1_85  = Y_ramRow[85];
  assign \U7/DATA1_86  = Y_ramRow[86];
  assign \U7/DATA1_87  = Y_ramRow[87];
  assign \U7/DATA1_88  = Y_ramRow[88];
  assign \U7/DATA1_89  = Y_ramRow[89];
  assign \U7/DATA1_90  = Y_ramRow[90];
  assign \U7/DATA1_91  = Y_ramRow[91];
  assign \U7/DATA1_92  = Y_ramRow[92];
  assign \U7/DATA1_93  = Y_ramRow[93];
  assign \U7/DATA1_94  = Y_ramRow[94];
  assign \U7/DATA1_95  = Y_ramRow[95];
  assign \U7/DATA1_96  = Y_ramRow[96];
  assign \U7/DATA1_97  = Y_ramRow[97];
  assign \U7/DATA1_98  = Y_ramRow[98];
  assign \U7/DATA1_99  = Y_ramRow[99];
  assign \U7/DATA1_100  = Y_ramRow[100];
  assign \U7/DATA1_101  = Y_ramRow[101];
  assign \U7/DATA1_102  = Y_ramRow[102];
  assign \U7/DATA1_103  = Y_ramRow[103];
  assign \U7/DATA1_104  = Y_ramRow[104];
  assign \U7/DATA1_105  = Y_ramRow[105];
  assign \U7/DATA1_106  = Y_ramRow[106];
  assign \U7/DATA1_107  = Y_ramRow[107];
  assign \U7/DATA1_108  = Y_ramRow[108];
  assign \U7/DATA1_109  = Y_ramRow[109];
  assign \U7/DATA1_110  = Y_ramRow[110];
  assign \U7/DATA1_111  = Y_ramRow[111];
  assign \U7/DATA1_128  = Y_ramRow[128];
  assign \U7/DATA1_129  = Y_ramRow[129];
  assign \U7/DATA1_130  = Y_ramRow[130];
  assign \U7/DATA1_131  = Y_ramRow[131];
  assign \U7/DATA1_132  = Y_ramRow[132];
  assign \U7/DATA1_133  = Y_ramRow[133];
  assign \U7/DATA1_134  = Y_ramRow[134];
  assign \U7/DATA1_135  = Y_ramRow[135];
  assign \U7/DATA1_136  = Y_ramRow[136];
  assign \U7/DATA1_137  = Y_ramRow[137];
  assign \U7/DATA1_138  = Y_ramRow[138];
  assign \U7/DATA1_139  = Y_ramRow[139];
  assign \U7/DATA1_140  = Y_ramRow[140];
  assign \U7/DATA1_141  = Y_ramRow[141];
  assign \U7/DATA1_142  = Y_ramRow[142];
  assign \U7/DATA1_143  = Y_ramRow[143];
  assign \U7/DATA1_144  = Y_ramRow[144];
  assign \U7/DATA1_145  = Y_ramRow[145];
  assign \U7/DATA1_146  = Y_ramRow[146];
  assign \U7/DATA1_147  = Y_ramRow[147];
  assign \U7/DATA1_148  = Y_ramRow[148];
  assign \U7/DATA1_149  = Y_ramRow[149];
  assign \U7/DATA1_150  = Y_ramRow[150];
  assign \U7/DATA1_151  = Y_ramRow[151];
  assign \U7/DATA1_152  = Y_ramRow[152];
  assign \U7/DATA1_153  = Y_ramRow[153];
  assign \U7/DATA1_154  = Y_ramRow[154];
  assign \U7/DATA1_155  = Y_ramRow[155];
  assign \U7/DATA1_156  = Y_ramRow[156];
  assign \U7/DATA1_157  = Y_ramRow[157];
  assign \U7/DATA1_158  = Y_ramRow[158];
  assign \U7/DATA1_159  = Y_ramRow[159];
  assign \U7/DATA1_160  = Y_ramRow[160];
  assign \U7/DATA1_161  = Y_ramRow[161];
  assign \U7/DATA1_162  = Y_ramRow[162];
  assign \U7/DATA1_163  = Y_ramRow[163];
  assign \U7/DATA1_164  = Y_ramRow[164];
  assign \U7/DATA1_165  = Y_ramRow[165];
  assign \U7/DATA1_166  = Y_ramRow[166];
  assign \U7/DATA1_167  = Y_ramRow[167];
  assign \U7/DATA1_168  = Y_ramRow[168];
  assign \U7/DATA1_169  = Y_ramRow[169];
  assign \U7/DATA1_170  = Y_ramRow[170];
  assign \U7/DATA1_171  = Y_ramRow[171];
  assign \U7/DATA1_172  = Y_ramRow[172];
  assign \U7/DATA1_173  = Y_ramRow[173];
  assign \U7/DATA1_174  = Y_ramRow[174];
  assign \U7/DATA1_175  = Y_ramRow[175];
  assign \U7/DATA1_192  = Element[0];
  assign \U7/DATA1_193  = Element[1];
  assign \U7/DATA1_194  = Element[2];
  assign \U7/DATA1_195  = Element[3];
  assign \U7/DATA1_196  = Element[4];
  assign \U7/DATA1_197  = Element[5];
  assign \U7/DATA1_198  = Element[6];
  assign \U7/DATA1_199  = Element[7];
  assign \U7/DATA1_200  = Element[8];
  assign \U7/DATA1_201  = Element[9];
  assign \U7/DATA1_202  = Element[10];
  assign \U7/DATA1_203  = Element[11];
  assign \U7/DATA1_204  = Element[12];
  assign \U7/DATA1_205  = Element[13];
  assign \U7/DATA1_206  = Element[14];
  assign \U7/DATA1_207  = Element[15];
  assign \U7/DATA1_208  = Element[16];
  assign \U7/DATA1_209  = Element[17];
  assign \U7/DATA1_210  = Element[18];
  assign \U7/DATA1_211  = Element[19];
  assign \U7/DATA1_212  = Element[20];
  assign \U7/DATA1_213  = Element[21];
  assign \U7/DATA1_214  = Element[22];
  assign \U7/DATA1_215  = Element[23];
  assign \U7/DATA1_216  = Element[24];
  assign \U7/DATA1_217  = Element[25];
  assign \U7/DATA1_218  = Element[26];
  assign \U7/DATA1_219  = Element[27];
  assign \U7/DATA1_220  = Element[28];
  assign \U7/DATA1_221  = Element[29];
  assign \U7/DATA1_222  = Element[30];
  assign \U7/DATA1_223  = Element[31];
  assign \U7/DATA1_224  = Element[32];
  assign \U7/DATA1_225  = Element[33];
  assign \U7/DATA1_226  = Element[34];
  assign \U7/DATA1_227  = Element[35];
  assign \U7/DATA1_228  = Element[36];
  assign \U7/DATA1_229  = Element[37];
  assign \U7/DATA1_230  = Element[38];
  assign \U7/DATA1_231  = Element[39];
  assign \U7/DATA1_232  = Element[40];
  assign \U7/DATA1_233  = Element[41];
  assign \U7/DATA1_234  = Element[42];
  assign \U7/DATA1_235  = Element[43];
  assign \U7/DATA1_236  = Element[44];
  assign \U7/DATA1_237  = Element[45];
  assign \U7/DATA1_238  = Element[46];
  assign \U7/DATA1_239  = Element[47];
  assign \U6/DATA1_192  = Y_ramRow[192];
  assign \U6/DATA1_193  = Y_ramRow[193];
  assign \U6/DATA1_194  = Y_ramRow[194];
  assign \U6/DATA1_195  = Y_ramRow[195];
  assign \U6/DATA1_196  = Y_ramRow[196];
  assign \U6/DATA1_197  = Y_ramRow[197];
  assign \U6/DATA1_198  = Y_ramRow[198];
  assign \U6/DATA1_199  = Y_ramRow[199];
  assign \U6/DATA1_200  = Y_ramRow[200];
  assign \U6/DATA1_201  = Y_ramRow[201];
  assign \U6/DATA1_202  = Y_ramRow[202];
  assign \U6/DATA1_203  = Y_ramRow[203];
  assign \U6/DATA1_204  = Y_ramRow[204];
  assign \U6/DATA1_205  = Y_ramRow[205];
  assign \U6/DATA1_206  = Y_ramRow[206];
  assign \U6/DATA1_207  = Y_ramRow[207];
  assign \U6/DATA1_208  = Y_ramRow[208];
  assign \U6/DATA1_209  = Y_ramRow[209];
  assign \U6/DATA1_210  = Y_ramRow[210];
  assign \U6/DATA1_211  = Y_ramRow[211];
  assign \U6/DATA1_212  = Y_ramRow[212];
  assign \U6/DATA1_213  = Y_ramRow[213];
  assign \U6/DATA1_214  = Y_ramRow[214];
  assign \U6/DATA1_215  = Y_ramRow[215];
  assign \U6/DATA1_216  = Y_ramRow[216];
  assign \U6/DATA1_217  = Y_ramRow[217];
  assign \U6/DATA1_218  = Y_ramRow[218];
  assign \U6/DATA1_219  = Y_ramRow[219];
  assign \U6/DATA1_220  = Y_ramRow[220];
  assign \U6/DATA1_221  = Y_ramRow[221];
  assign \U6/DATA1_222  = Y_ramRow[222];
  assign \U6/DATA1_223  = Y_ramRow[223];
  assign \U6/DATA1_224  = Y_ramRow[224];
  assign \U6/DATA1_225  = Y_ramRow[225];
  assign \U6/DATA1_226  = Y_ramRow[226];
  assign \U6/DATA1_227  = Y_ramRow[227];
  assign \U6/DATA1_228  = Y_ramRow[228];
  assign \U6/DATA1_229  = Y_ramRow[229];
  assign \U6/DATA1_230  = Y_ramRow[230];
  assign \U6/DATA1_231  = Y_ramRow[231];
  assign \U6/DATA1_232  = Y_ramRow[232];
  assign \U6/DATA1_233  = Y_ramRow[233];
  assign \U6/DATA1_234  = Y_ramRow[234];
  assign \U6/DATA1_235  = Y_ramRow[235];
  assign \U6/DATA1_236  = Y_ramRow[236];
  assign \U6/DATA1_237  = Y_ramRow[237];
  assign \U6/DATA1_238  = Y_ramRow[238];
  assign \U6/DATA1_239  = Y_ramRow[239];
  assign PaddedRow[0] = \U4/Z_0 ;
  assign PaddedRow[1] = \U4/Z_1 ;
  assign PaddedRow[2] = \U4/Z_2 ;
  assign PaddedRow[3] = \U4/Z_3 ;
  assign PaddedRow[4] = \U4/Z_4 ;
  assign PaddedRow[5] = \U4/Z_5 ;
  assign PaddedRow[6] = \U4/Z_6 ;
  assign PaddedRow[7] = \U4/Z_7 ;
  assign PaddedRow[8] = \U4/Z_8 ;
  assign PaddedRow[9] = \U4/Z_9 ;
  assign PaddedRow[10] = \U4/Z_10 ;
  assign PaddedRow[11] = \U4/Z_11 ;
  assign PaddedRow[12] = \U4/Z_12 ;
  assign PaddedRow[13] = \U4/Z_13 ;
  assign PaddedRow[14] = \U4/Z_14 ;
  assign PaddedRow[15] = \U4/Z_15 ;
  assign PaddedRow[16] = \U4/Z_16 ;
  assign PaddedRow[17] = \U4/Z_17 ;
  assign PaddedRow[18] = \U4/Z_18 ;
  assign PaddedRow[19] = \U4/Z_19 ;
  assign PaddedRow[20] = \U4/Z_20 ;
  assign PaddedRow[21] = \U4/Z_21 ;
  assign PaddedRow[22] = \U4/Z_22 ;
  assign PaddedRow[23] = \U4/Z_23 ;
  assign PaddedRow[24] = \U4/Z_24 ;
  assign PaddedRow[25] = \U4/Z_25 ;
  assign PaddedRow[26] = \U4/Z_26 ;
  assign PaddedRow[27] = \U4/Z_27 ;
  assign PaddedRow[28] = \U4/Z_28 ;
  assign PaddedRow[29] = \U4/Z_29 ;
  assign PaddedRow[30] = \U4/Z_30 ;
  assign PaddedRow[31] = \U4/Z_31 ;
  assign PaddedRow[32] = \U4/Z_32 ;
  assign PaddedRow[33] = \U4/Z_33 ;
  assign PaddedRow[34] = \U4/Z_34 ;
  assign PaddedRow[35] = \U4/Z_35 ;
  assign PaddedRow[36] = \U4/Z_36 ;
  assign PaddedRow[37] = \U4/Z_37 ;
  assign PaddedRow[38] = \U4/Z_38 ;
  assign PaddedRow[39] = \U4/Z_39 ;
  assign PaddedRow[40] = \U4/Z_40 ;
  assign PaddedRow[41] = \U4/Z_41 ;
  assign PaddedRow[42] = \U4/Z_42 ;
  assign PaddedRow[43] = \U4/Z_43 ;
  assign PaddedRow[44] = \U4/Z_44 ;
  assign PaddedRow[45] = \U4/Z_45 ;
  assign PaddedRow[46] = \U4/Z_46 ;
  assign PaddedRow[47] = \U4/Z_47 ;
  assign \U4/Z_48  = Y_ramRow[48];
  assign \U4/Z_49  = Y_ramRow[49];
  assign \U4/Z_50  = Y_ramRow[50];
  assign \U4/Z_51  = Y_ramRow[51];
  assign \U4/Z_52  = Y_ramRow[52];
  assign \U4/Z_53  = Y_ramRow[53];
  assign \U4/Z_54  = Y_ramRow[54];
  assign \U4/Z_55  = Y_ramRow[55];
  assign \U4/Z_56  = Y_ramRow[56];
  assign \U4/Z_57  = Y_ramRow[57];
  assign \U4/Z_58  = Y_ramRow[58];
  assign \U4/Z_59  = Y_ramRow[59];
  assign \U4/Z_60  = Y_ramRow[60];
  assign \U4/Z_61  = Y_ramRow[61];
  assign \U4/Z_62  = Y_ramRow[62];
  assign \U4/Z_63  = Y_ramRow[63];
  assign PaddedRow[64] = \U4/Z_64 ;
  assign PaddedRow[65] = \U4/Z_65 ;
  assign PaddedRow[66] = \U4/Z_66 ;
  assign PaddedRow[67] = \U4/Z_67 ;
  assign PaddedRow[68] = \U4/Z_68 ;
  assign PaddedRow[69] = \U4/Z_69 ;
  assign PaddedRow[70] = \U4/Z_70 ;
  assign PaddedRow[71] = \U4/Z_71 ;
  assign PaddedRow[72] = \U4/Z_72 ;
  assign PaddedRow[73] = \U4/Z_73 ;
  assign PaddedRow[74] = \U4/Z_74 ;
  assign PaddedRow[75] = \U4/Z_75 ;
  assign PaddedRow[76] = \U4/Z_76 ;
  assign PaddedRow[77] = \U4/Z_77 ;
  assign PaddedRow[78] = \U4/Z_78 ;
  assign PaddedRow[79] = \U4/Z_79 ;
  assign PaddedRow[80] = \U4/Z_80 ;
  assign PaddedRow[81] = \U4/Z_81 ;
  assign PaddedRow[82] = \U4/Z_82 ;
  assign PaddedRow[83] = \U4/Z_83 ;
  assign PaddedRow[84] = \U4/Z_84 ;
  assign PaddedRow[85] = \U4/Z_85 ;
  assign PaddedRow[86] = \U4/Z_86 ;
  assign PaddedRow[87] = \U4/Z_87 ;
  assign PaddedRow[88] = \U4/Z_88 ;
  assign PaddedRow[89] = \U4/Z_89 ;
  assign PaddedRow[90] = \U4/Z_90 ;
  assign PaddedRow[91] = \U4/Z_91 ;
  assign PaddedRow[92] = \U4/Z_92 ;
  assign PaddedRow[93] = \U4/Z_93 ;
  assign PaddedRow[94] = \U4/Z_94 ;
  assign PaddedRow[95] = \U4/Z_95 ;
  assign PaddedRow[96] = \U4/Z_96 ;
  assign PaddedRow[97] = \U4/Z_97 ;
  assign PaddedRow[98] = \U4/Z_98 ;
  assign PaddedRow[99] = \U4/Z_99 ;
  assign PaddedRow[100] = \U4/Z_100 ;
  assign PaddedRow[101] = \U4/Z_101 ;
  assign PaddedRow[102] = \U4/Z_102 ;
  assign PaddedRow[103] = \U4/Z_103 ;
  assign PaddedRow[104] = \U4/Z_104 ;
  assign PaddedRow[105] = \U4/Z_105 ;
  assign PaddedRow[106] = \U4/Z_106 ;
  assign PaddedRow[107] = \U4/Z_107 ;
  assign PaddedRow[108] = \U4/Z_108 ;
  assign PaddedRow[109] = \U4/Z_109 ;
  assign PaddedRow[110] = \U4/Z_110 ;
  assign PaddedRow[111] = \U4/Z_111 ;
  assign \U4/Z_112  = Y_ramRow[112];
  assign \U4/Z_113  = Y_ramRow[113];
  assign \U4/Z_114  = Y_ramRow[114];
  assign \U4/Z_115  = Y_ramRow[115];
  assign \U4/Z_116  = Y_ramRow[116];
  assign \U4/Z_117  = Y_ramRow[117];
  assign \U4/Z_118  = Y_ramRow[118];
  assign \U4/Z_119  = Y_ramRow[119];
  assign \U4/Z_120  = Y_ramRow[120];
  assign \U4/Z_121  = Y_ramRow[121];
  assign \U4/Z_122  = Y_ramRow[122];
  assign \U4/Z_123  = Y_ramRow[123];
  assign \U4/Z_124  = Y_ramRow[124];
  assign \U4/Z_125  = Y_ramRow[125];
  assign \U4/Z_126  = Y_ramRow[126];
  assign \U4/Z_127  = Y_ramRow[127];
  assign PaddedRow[128] = \U4/Z_128 ;
  assign PaddedRow[129] = \U4/Z_129 ;
  assign PaddedRow[130] = \U4/Z_130 ;
  assign PaddedRow[131] = \U4/Z_131 ;
  assign PaddedRow[132] = \U4/Z_132 ;
  assign PaddedRow[133] = \U4/Z_133 ;
  assign PaddedRow[134] = \U4/Z_134 ;
  assign PaddedRow[135] = \U4/Z_135 ;
  assign PaddedRow[136] = \U4/Z_136 ;
  assign PaddedRow[137] = \U4/Z_137 ;
  assign PaddedRow[138] = \U4/Z_138 ;
  assign PaddedRow[139] = \U4/Z_139 ;
  assign PaddedRow[140] = \U4/Z_140 ;
  assign PaddedRow[141] = \U4/Z_141 ;
  assign PaddedRow[142] = \U4/Z_142 ;
  assign PaddedRow[143] = \U4/Z_143 ;
  assign PaddedRow[144] = \U4/Z_144 ;
  assign PaddedRow[145] = \U4/Z_145 ;
  assign PaddedRow[146] = \U4/Z_146 ;
  assign PaddedRow[147] = \U4/Z_147 ;
  assign PaddedRow[148] = \U4/Z_148 ;
  assign PaddedRow[149] = \U4/Z_149 ;
  assign PaddedRow[150] = \U4/Z_150 ;
  assign PaddedRow[151] = \U4/Z_151 ;
  assign PaddedRow[152] = \U4/Z_152 ;
  assign PaddedRow[153] = \U4/Z_153 ;
  assign PaddedRow[154] = \U4/Z_154 ;
  assign PaddedRow[155] = \U4/Z_155 ;
  assign PaddedRow[156] = \U4/Z_156 ;
  assign PaddedRow[157] = \U4/Z_157 ;
  assign PaddedRow[158] = \U4/Z_158 ;
  assign PaddedRow[159] = \U4/Z_159 ;
  assign PaddedRow[160] = \U4/Z_160 ;
  assign PaddedRow[161] = \U4/Z_161 ;
  assign PaddedRow[162] = \U4/Z_162 ;
  assign PaddedRow[163] = \U4/Z_163 ;
  assign PaddedRow[164] = \U4/Z_164 ;
  assign PaddedRow[165] = \U4/Z_165 ;
  assign PaddedRow[166] = \U4/Z_166 ;
  assign PaddedRow[167] = \U4/Z_167 ;
  assign PaddedRow[168] = \U4/Z_168 ;
  assign PaddedRow[169] = \U4/Z_169 ;
  assign PaddedRow[170] = \U4/Z_170 ;
  assign PaddedRow[171] = \U4/Z_171 ;
  assign PaddedRow[172] = \U4/Z_172 ;
  assign PaddedRow[173] = \U4/Z_173 ;
  assign PaddedRow[174] = \U4/Z_174 ;
  assign PaddedRow[175] = \U4/Z_175 ;
  assign \U4/Z_176  = Y_ramRow[176];
  assign \U4/Z_177  = Y_ramRow[177];
  assign \U4/Z_178  = Y_ramRow[178];
  assign \U4/Z_179  = Y_ramRow[179];
  assign \U4/Z_180  = Y_ramRow[180];
  assign \U4/Z_181  = Y_ramRow[181];
  assign \U4/Z_182  = Y_ramRow[182];
  assign \U4/Z_183  = Y_ramRow[183];
  assign \U4/Z_184  = Y_ramRow[184];
  assign \U4/Z_185  = Y_ramRow[185];
  assign \U4/Z_186  = Y_ramRow[186];
  assign \U4/Z_187  = Y_ramRow[187];
  assign \U4/Z_188  = Y_ramRow[188];
  assign \U4/Z_189  = Y_ramRow[189];
  assign \U4/Z_190  = Y_ramRow[190];
  assign \U4/Z_191  = Y_ramRow[191];
  assign PaddedRow[192] = \U4/Z_192 ;
  assign PaddedRow[193] = \U4/Z_193 ;
  assign PaddedRow[194] = \U4/Z_194 ;
  assign PaddedRow[195] = \U4/Z_195 ;
  assign PaddedRow[196] = \U4/Z_196 ;
  assign PaddedRow[197] = \U4/Z_197 ;
  assign PaddedRow[198] = \U4/Z_198 ;
  assign PaddedRow[199] = \U4/Z_199 ;
  assign PaddedRow[200] = \U4/Z_200 ;
  assign PaddedRow[201] = \U4/Z_201 ;
  assign PaddedRow[202] = \U4/Z_202 ;
  assign PaddedRow[203] = \U4/Z_203 ;
  assign PaddedRow[204] = \U4/Z_204 ;
  assign PaddedRow[205] = \U4/Z_205 ;
  assign PaddedRow[206] = \U4/Z_206 ;
  assign PaddedRow[207] = \U4/Z_207 ;
  assign PaddedRow[208] = \U4/Z_208 ;
  assign PaddedRow[209] = \U4/Z_209 ;
  assign PaddedRow[210] = \U4/Z_210 ;
  assign PaddedRow[211] = \U4/Z_211 ;
  assign PaddedRow[212] = \U4/Z_212 ;
  assign PaddedRow[213] = \U4/Z_213 ;
  assign PaddedRow[214] = \U4/Z_214 ;
  assign PaddedRow[215] = \U4/Z_215 ;
  assign PaddedRow[216] = \U4/Z_216 ;
  assign PaddedRow[217] = \U4/Z_217 ;
  assign PaddedRow[218] = \U4/Z_218 ;
  assign PaddedRow[219] = \U4/Z_219 ;
  assign PaddedRow[220] = \U4/Z_220 ;
  assign PaddedRow[221] = \U4/Z_221 ;
  assign PaddedRow[222] = \U4/Z_222 ;
  assign PaddedRow[223] = \U4/Z_223 ;
  assign PaddedRow[224] = \U4/Z_224 ;
  assign PaddedRow[225] = \U4/Z_225 ;
  assign PaddedRow[226] = \U4/Z_226 ;
  assign PaddedRow[227] = \U4/Z_227 ;
  assign PaddedRow[228] = \U4/Z_228 ;
  assign PaddedRow[229] = \U4/Z_229 ;
  assign PaddedRow[230] = \U4/Z_230 ;
  assign PaddedRow[231] = \U4/Z_231 ;
  assign PaddedRow[232] = \U4/Z_232 ;
  assign PaddedRow[233] = \U4/Z_233 ;
  assign PaddedRow[234] = \U4/Z_234 ;
  assign PaddedRow[235] = \U4/Z_235 ;
  assign PaddedRow[236] = \U4/Z_236 ;
  assign PaddedRow[237] = \U4/Z_237 ;
  assign PaddedRow[238] = \U4/Z_238 ;
  assign PaddedRow[239] = \U4/Z_239 ;
  assign \U4/Z_240  = Y_ramRow[240];
  assign \U4/Z_241  = Y_ramRow[241];
  assign \U4/Z_242  = Y_ramRow[242];
  assign \U4/Z_243  = Y_ramRow[243];
  assign \U4/Z_244  = Y_ramRow[244];
  assign \U4/Z_245  = Y_ramRow[245];
  assign \U4/Z_246  = Y_ramRow[246];
  assign \U4/Z_247  = Y_ramRow[247];
  assign \U4/Z_248  = Y_ramRow[248];
  assign \U4/Z_249  = Y_ramRow[249];
  assign \U4/Z_250  = Y_ramRow[250];
  assign \U4/Z_251  = Y_ramRow[251];
  assign \U4/Z_252  = Y_ramRow[252];
  assign \U4/Z_253  = Y_ramRow[253];
  assign \U4/Z_254  = Y_ramRow[254];
  assign \U4/Z_255  = Y_ramRow[255];

  NAND2_X2 U4 ( .A1(\U7/DATA1_99 ), .A2(n1363), .ZN(n51) );
  NAND2_X2 U6 ( .A1(\U7/DATA1_98 ), .A2(n1363), .ZN(n53) );
  NAND2_X2 U8 ( .A1(\U7/DATA1_97 ), .A2(n1363), .ZN(n54) );
  NAND2_X2 U10 ( .A1(\U7/DATA1_96 ), .A2(n1363), .ZN(n55) );
  NAND2_X2 U12 ( .A1(\U7/DATA1_95 ), .A2(n1363), .ZN(n56) );
  NAND2_X2 U14 ( .A1(\U7/DATA1_94 ), .A2(n1363), .ZN(n57) );
  NAND2_X2 U16 ( .A1(\U7/DATA1_93 ), .A2(n1363), .ZN(n58) );
  NAND2_X2 U18 ( .A1(\U7/DATA1_92 ), .A2(n1363), .ZN(n59) );
  NAND2_X2 U20 ( .A1(\U7/DATA1_91 ), .A2(n1363), .ZN(n60) );
  NAND2_X2 U22 ( .A1(\U7/DATA1_90 ), .A2(n1363), .ZN(n61) );
  NAND2_X2 U24 ( .A1(\U7/DATA1_9 ), .A2(n1364), .ZN(n63) );
  NAND2_X2 U26 ( .A1(\U7/DATA1_89 ), .A2(n1363), .ZN(n65) );
  NAND2_X2 U28 ( .A1(\U7/DATA1_88 ), .A2(n1363), .ZN(n66) );
  NAND2_X2 U30 ( .A1(\U7/DATA1_87 ), .A2(n1363), .ZN(n67) );
  NAND2_X2 U32 ( .A1(\U7/DATA1_86 ), .A2(n1363), .ZN(n68) );
  NAND2_X2 U34 ( .A1(\U7/DATA1_85 ), .A2(n1363), .ZN(n69) );
  NAND2_X2 U36 ( .A1(\U7/DATA1_84 ), .A2(n1363), .ZN(n70) );
  NAND2_X2 U38 ( .A1(\U7/DATA1_83 ), .A2(n1363), .ZN(n71) );
  NAND2_X2 U40 ( .A1(\U7/DATA1_82 ), .A2(n1363), .ZN(n72) );
  NAND2_X2 U42 ( .A1(\U7/DATA1_81 ), .A2(n1363), .ZN(n73) );
  NAND2_X2 U44 ( .A1(\U7/DATA1_80 ), .A2(n1363), .ZN(n74) );
  NAND2_X2 U46 ( .A1(\U7/DATA1_8 ), .A2(n1364), .ZN(n75) );
  NAND2_X2 U48 ( .A1(\U7/DATA1_79 ), .A2(n1363), .ZN(n76) );
  NAND2_X2 U50 ( .A1(\U7/DATA1_78 ), .A2(n1363), .ZN(n77) );
  NAND2_X2 U52 ( .A1(\U7/DATA1_77 ), .A2(n1363), .ZN(n78) );
  NAND2_X2 U54 ( .A1(\U7/DATA1_76 ), .A2(n1363), .ZN(n79) );
  NAND2_X2 U56 ( .A1(\U7/DATA1_75 ), .A2(n1363), .ZN(n80) );
  NAND2_X2 U58 ( .A1(\U7/DATA1_74 ), .A2(n1363), .ZN(n81) );
  NAND2_X2 U60 ( .A1(\U7/DATA1_73 ), .A2(n1363), .ZN(n82) );
  NAND2_X2 U62 ( .A1(\U7/DATA1_72 ), .A2(n1363), .ZN(n83) );
  NAND2_X2 U64 ( .A1(\U7/DATA1_71 ), .A2(n1363), .ZN(n84) );
  NAND2_X2 U66 ( .A1(\U7/DATA1_70 ), .A2(n1363), .ZN(n85) );
  NAND2_X2 U68 ( .A1(\U7/DATA1_7 ), .A2(n1364), .ZN(n86) );
  NAND2_X2 U70 ( .A1(\U7/DATA1_69 ), .A2(n1363), .ZN(n87) );
  NAND2_X2 U72 ( .A1(\U7/DATA1_68 ), .A2(n1363), .ZN(n88) );
  NAND2_X2 U74 ( .A1(\U7/DATA1_67 ), .A2(n1363), .ZN(n89) );
  NAND2_X2 U76 ( .A1(\U7/DATA1_66 ), .A2(n1363), .ZN(n90) );
  NAND2_X2 U78 ( .A1(\U7/DATA1_65 ), .A2(n1363), .ZN(n91) );
  NAND2_X2 U80 ( .A1(\U7/DATA1_64 ), .A2(n1363), .ZN(n92) );
  NAND2_X2 U82 ( .A1(\U7/DATA1_6 ), .A2(n1364), .ZN(n93) );
  NAND2_X2 U84 ( .A1(\U7/DATA1_5 ), .A2(n1364), .ZN(n94) );
  NAND2_X2 U86 ( .A1(\U7/DATA1_47 ), .A2(n1364), .ZN(n95) );
  NAND2_X2 U88 ( .A1(\U7/DATA1_46 ), .A2(n1364), .ZN(n96) );
  NAND2_X2 U90 ( .A1(\U7/DATA1_45 ), .A2(n1364), .ZN(n97) );
  NAND2_X2 U92 ( .A1(\U7/DATA1_44 ), .A2(n1364), .ZN(n98) );
  NAND2_X2 U94 ( .A1(\U7/DATA1_43 ), .A2(n1364), .ZN(n99) );
  NAND2_X2 U96 ( .A1(\U7/DATA1_42 ), .A2(n1364), .ZN(n100) );
  NAND2_X2 U98 ( .A1(\U7/DATA1_41 ), .A2(n1364), .ZN(n101) );
  NAND2_X2 U100 ( .A1(\U7/DATA1_40 ), .A2(n1364), .ZN(n102) );
  NAND2_X2 U102 ( .A1(\U7/DATA1_4 ), .A2(n1364), .ZN(n103) );
  NAND2_X2 U104 ( .A1(\U7/DATA1_39 ), .A2(n1364), .ZN(n104) );
  NAND2_X2 U106 ( .A1(\U7/DATA1_38 ), .A2(n1364), .ZN(n105) );
  NAND2_X2 U108 ( .A1(\U7/DATA1_37 ), .A2(n1364), .ZN(n106) );
  NAND2_X2 U110 ( .A1(\U7/DATA1_36 ), .A2(n1364), .ZN(n107) );
  NAND2_X2 U112 ( .A1(\U7/DATA1_35 ), .A2(n1364), .ZN(n108) );
  NAND2_X2 U114 ( .A1(\U7/DATA1_34 ), .A2(n1364), .ZN(n109) );
  NAND2_X2 U116 ( .A1(\U7/DATA1_33 ), .A2(n1364), .ZN(n110) );
  NAND2_X2 U118 ( .A1(\U7/DATA1_32 ), .A2(n1364), .ZN(n111) );
  NAND2_X2 U120 ( .A1(\U7/DATA1_31 ), .A2(n1364), .ZN(n112) );
  NAND2_X2 U122 ( .A1(\U7/DATA1_30 ), .A2(n1364), .ZN(n113) );
  NAND2_X2 U124 ( .A1(\U7/DATA1_3 ), .A2(n1364), .ZN(n114) );
  NAND2_X2 U126 ( .A1(\U7/DATA1_29 ), .A2(n1364), .ZN(n115) );
  NAND2_X2 U128 ( .A1(\U7/DATA1_28 ), .A2(n1364), .ZN(n116) );
  NAND2_X2 U130 ( .A1(\U7/DATA1_27 ), .A2(n1364), .ZN(n117) );
  NAND2_X2 U132 ( .A1(\U7/DATA1_26 ), .A2(n1364), .ZN(n118) );
  NAND2_X2 U134 ( .A1(\U7/DATA1_25 ), .A2(n1364), .ZN(n119) );
  NAND2_X2 U136 ( .A1(\U7/DATA1_24 ), .A2(n1364), .ZN(n120) );
  NAND2_X2 U138 ( .A1(\U6/DATA1_239 ), .A2(n1433), .ZN(n122) );
  NAND2_X2 U140 ( .A1(\U6/DATA1_238 ), .A2(n1434), .ZN(n123) );
  NAND2_X2 U142 ( .A1(\U6/DATA1_237 ), .A2(n1434), .ZN(n124) );
  NAND2_X2 U144 ( .A1(\U6/DATA1_236 ), .A2(n1434), .ZN(n125) );
  NAND2_X2 U146 ( .A1(\U6/DATA1_235 ), .A2(n1434), .ZN(n126) );
  NAND2_X2 U148 ( .A1(\U6/DATA1_234 ), .A2(n1434), .ZN(n127) );
  NAND2_X2 U150 ( .A1(\U6/DATA1_233 ), .A2(n1434), .ZN(n128) );
  NAND2_X2 U152 ( .A1(\U6/DATA1_232 ), .A2(n1433), .ZN(n129) );
  NAND2_X2 U154 ( .A1(\U6/DATA1_231 ), .A2(n1434), .ZN(n130) );
  NAND2_X2 U156 ( .A1(\U6/DATA1_230 ), .A2(n1434), .ZN(n131) );
  NAND2_X2 U158 ( .A1(\U7/DATA1_23 ), .A2(n1364), .ZN(n132) );
  NAND2_X2 U160 ( .A1(\U6/DATA1_229 ), .A2(n1434), .ZN(n133) );
  NAND2_X2 U162 ( .A1(\U6/DATA1_228 ), .A2(n1434), .ZN(n134) );
  NAND2_X2 U164 ( .A1(\U6/DATA1_227 ), .A2(n1434), .ZN(n135) );
  NAND2_X2 U166 ( .A1(\U6/DATA1_226 ), .A2(n1434), .ZN(n136) );
  NAND2_X2 U168 ( .A1(\U6/DATA1_225 ), .A2(n1434), .ZN(n137) );
  NAND2_X2 U170 ( .A1(\U6/DATA1_224 ), .A2(n1434), .ZN(n138) );
  NAND2_X2 U172 ( .A1(\U6/DATA1_223 ), .A2(n1434), .ZN(n139) );
  NAND2_X2 U174 ( .A1(\U6/DATA1_222 ), .A2(n1434), .ZN(n140) );
  NAND2_X2 U176 ( .A1(\U6/DATA1_221 ), .A2(n1434), .ZN(n141) );
  NAND2_X2 U178 ( .A1(\U6/DATA1_220 ), .A2(n1434), .ZN(n142) );
  NAND2_X2 U180 ( .A1(\U7/DATA1_22 ), .A2(n1364), .ZN(n143) );
  NAND2_X2 U182 ( .A1(\U6/DATA1_219 ), .A2(n1434), .ZN(n144) );
  NAND2_X2 U184 ( .A1(\U6/DATA1_218 ), .A2(n1434), .ZN(n145) );
  NAND2_X2 U186 ( .A1(\U6/DATA1_217 ), .A2(n1434), .ZN(n146) );
  NAND2_X2 U188 ( .A1(\U6/DATA1_216 ), .A2(n1434), .ZN(n147) );
  NAND2_X2 U190 ( .A1(\U6/DATA1_215 ), .A2(n1434), .ZN(n148) );
  NAND2_X2 U192 ( .A1(\U6/DATA1_214 ), .A2(n1434), .ZN(n149) );
  NAND2_X2 U194 ( .A1(\U6/DATA1_213 ), .A2(n1434), .ZN(n150) );
  NAND2_X2 U196 ( .A1(\U6/DATA1_212 ), .A2(n1434), .ZN(n151) );
  NAND2_X2 U198 ( .A1(\U6/DATA1_211 ), .A2(n1434), .ZN(n152) );
  NAND2_X2 U200 ( .A1(\U6/DATA1_210 ), .A2(n1434), .ZN(n153) );
  NAND2_X2 U202 ( .A1(\U7/DATA1_21 ), .A2(n1364), .ZN(n154) );
  NAND2_X2 U204 ( .A1(\U6/DATA1_209 ), .A2(n1434), .ZN(n155) );
  NAND2_X2 U206 ( .A1(\U6/DATA1_208 ), .A2(n1434), .ZN(n156) );
  NAND2_X2 U208 ( .A1(\U6/DATA1_207 ), .A2(n1434), .ZN(n157) );
  NAND2_X2 U210 ( .A1(\U6/DATA1_206 ), .A2(n1434), .ZN(n158) );
  NAND2_X2 U212 ( .A1(\U6/DATA1_205 ), .A2(n1434), .ZN(n159) );
  NAND2_X2 U214 ( .A1(\U6/DATA1_204 ), .A2(n1434), .ZN(n160) );
  NAND2_X2 U216 ( .A1(\U6/DATA1_203 ), .A2(n1434), .ZN(n161) );
  NAND2_X2 U218 ( .A1(\U6/DATA1_202 ), .A2(n1434), .ZN(n162) );
  NAND2_X2 U220 ( .A1(\U6/DATA1_201 ), .A2(n1434), .ZN(n163) );
  NAND2_X2 U222 ( .A1(\U6/DATA1_200 ), .A2(n1434), .ZN(n164) );
  NAND2_X2 U224 ( .A1(\U7/DATA1_20 ), .A2(n1364), .ZN(n165) );
  NAND2_X2 U226 ( .A1(\U7/DATA1_2 ), .A2(n1364), .ZN(n166) );
  NAND2_X2 U228 ( .A1(\U6/DATA1_199 ), .A2(n1434), .ZN(n167) );
  NAND2_X2 U230 ( .A1(\U6/DATA1_198 ), .A2(n1434), .ZN(n168) );
  NAND2_X2 U232 ( .A1(\U6/DATA1_197 ), .A2(n1434), .ZN(n169) );
  NAND2_X2 U234 ( .A1(\U6/DATA1_196 ), .A2(n1434), .ZN(n170) );
  NAND2_X2 U236 ( .A1(\U6/DATA1_195 ), .A2(n1434), .ZN(n171) );
  NAND2_X2 U238 ( .A1(\U6/DATA1_194 ), .A2(n1434), .ZN(n172) );
  NAND2_X2 U240 ( .A1(\U6/DATA1_193 ), .A2(n1434), .ZN(n173) );
  NAND2_X2 U242 ( .A1(\U6/DATA1_192 ), .A2(n1434), .ZN(n174) );
  NAND2_X2 U245 ( .A1(\U7/DATA1_19 ), .A2(n1364), .ZN(n176) );
  NAND2_X2 U247 ( .A1(\U7/DATA1_18 ), .A2(n1364), .ZN(n177) );
  NAND2_X2 U249 ( .A1(\U7/DATA1_175 ), .A2(n1432), .ZN(n178) );
  NAND2_X2 U251 ( .A1(\U7/DATA1_174 ), .A2(n1432), .ZN(n179) );
  NAND2_X2 U253 ( .A1(\U7/DATA1_173 ), .A2(n1432), .ZN(n180) );
  NAND2_X2 U255 ( .A1(\U7/DATA1_172 ), .A2(n1432), .ZN(n181) );
  NAND2_X2 U257 ( .A1(\U7/DATA1_171 ), .A2(n1432), .ZN(n182) );
  NAND2_X2 U259 ( .A1(\U7/DATA1_170 ), .A2(n1432), .ZN(n183) );
  NAND2_X2 U261 ( .A1(\U7/DATA1_17 ), .A2(n1364), .ZN(n184) );
  NAND2_X2 U263 ( .A1(\U7/DATA1_169 ), .A2(n1432), .ZN(n185) );
  NAND2_X2 U265 ( .A1(\U7/DATA1_168 ), .A2(n1432), .ZN(n186) );
  NAND2_X2 U267 ( .A1(\U7/DATA1_167 ), .A2(n1432), .ZN(n187) );
  NAND2_X2 U269 ( .A1(\U7/DATA1_166 ), .A2(n1432), .ZN(n188) );
  NAND2_X2 U271 ( .A1(\U7/DATA1_165 ), .A2(n1432), .ZN(n189) );
  NAND2_X2 U273 ( .A1(\U7/DATA1_164 ), .A2(n1432), .ZN(n190) );
  NAND2_X2 U275 ( .A1(\U7/DATA1_163 ), .A2(n1432), .ZN(n191) );
  NAND2_X2 U277 ( .A1(\U7/DATA1_162 ), .A2(n1432), .ZN(n192) );
  NAND2_X2 U279 ( .A1(\U7/DATA1_161 ), .A2(n1432), .ZN(n193) );
  NAND2_X2 U281 ( .A1(\U7/DATA1_160 ), .A2(n1432), .ZN(n194) );
  NAND2_X2 U283 ( .A1(\U7/DATA1_16 ), .A2(n1364), .ZN(n195) );
  NAND2_X2 U285 ( .A1(\U7/DATA1_159 ), .A2(n1432), .ZN(n196) );
  NAND2_X2 U287 ( .A1(\U7/DATA1_158 ), .A2(n1432), .ZN(n197) );
  NAND2_X2 U289 ( .A1(\U7/DATA1_157 ), .A2(n1432), .ZN(n198) );
  NAND2_X2 U291 ( .A1(\U7/DATA1_156 ), .A2(n1432), .ZN(n199) );
  NAND2_X2 U293 ( .A1(\U7/DATA1_155 ), .A2(n1432), .ZN(n200) );
  NAND2_X2 U295 ( .A1(\U7/DATA1_154 ), .A2(n1432), .ZN(n201) );
  NAND2_X2 U297 ( .A1(\U7/DATA1_153 ), .A2(n1432), .ZN(n202) );
  NAND2_X2 U299 ( .A1(\U7/DATA1_152 ), .A2(n1432), .ZN(n203) );
  NAND2_X2 U301 ( .A1(\U7/DATA1_151 ), .A2(n1432), .ZN(n204) );
  NAND2_X2 U303 ( .A1(\U7/DATA1_150 ), .A2(n1432), .ZN(n205) );
  NAND2_X2 U305 ( .A1(\U7/DATA1_15 ), .A2(n1364), .ZN(n206) );
  NAND2_X2 U307 ( .A1(\U7/DATA1_149 ), .A2(n1432), .ZN(n207) );
  NAND2_X2 U309 ( .A1(\U7/DATA1_148 ), .A2(n175), .ZN(n208) );
  NAND2_X2 U311 ( .A1(\U7/DATA1_147 ), .A2(n175), .ZN(n209) );
  NAND2_X2 U313 ( .A1(\U7/DATA1_146 ), .A2(n175), .ZN(n210) );
  NAND2_X2 U315 ( .A1(\U7/DATA1_145 ), .A2(n175), .ZN(n211) );
  NAND2_X2 U317 ( .A1(\U7/DATA1_144 ), .A2(n175), .ZN(n212) );
  NAND2_X2 U319 ( .A1(\U7/DATA1_143 ), .A2(n175), .ZN(n213) );
  NAND2_X2 U321 ( .A1(\U7/DATA1_142 ), .A2(n175), .ZN(n214) );
  NAND2_X2 U323 ( .A1(\U7/DATA1_141 ), .A2(n175), .ZN(n215) );
  NAND2_X2 U325 ( .A1(\U7/DATA1_140 ), .A2(n175), .ZN(n216) );
  NAND2_X2 U327 ( .A1(\U7/DATA1_14 ), .A2(n1364), .ZN(n217) );
  NAND2_X2 U329 ( .A1(\U7/DATA1_139 ), .A2(n175), .ZN(n218) );
  NAND2_X2 U331 ( .A1(\U7/DATA1_138 ), .A2(n175), .ZN(n219) );
  NAND2_X2 U333 ( .A1(\U7/DATA1_137 ), .A2(n175), .ZN(n220) );
  NAND2_X2 U335 ( .A1(\U7/DATA1_136 ), .A2(n175), .ZN(n221) );
  NAND2_X2 U337 ( .A1(\U7/DATA1_135 ), .A2(n1432), .ZN(n222) );
  NAND2_X2 U339 ( .A1(\U7/DATA1_134 ), .A2(n1432), .ZN(n223) );
  NAND2_X2 U341 ( .A1(\U7/DATA1_133 ), .A2(n1432), .ZN(n224) );
  NAND2_X2 U343 ( .A1(\U7/DATA1_132 ), .A2(n1431), .ZN(n225) );
  NAND2_X2 U345 ( .A1(\U7/DATA1_131 ), .A2(n1431), .ZN(n226) );
  NAND2_X2 U347 ( .A1(\U7/DATA1_130 ), .A2(n1431), .ZN(n227) );
  NAND2_X2 U349 ( .A1(\U7/DATA1_13 ), .A2(n1364), .ZN(n228) );
  NAND2_X2 U351 ( .A1(\U7/DATA1_129 ), .A2(n1431), .ZN(n229) );
  NAND2_X2 U353 ( .A1(\U7/DATA1_128 ), .A2(n1432), .ZN(n230) );
  NAND2_X2 U354 ( .A1(PosElement[0]), .A2(n1485), .ZN(n175) );
  NAND2_X2 U356 ( .A1(\U7/DATA1_12 ), .A2(n1364), .ZN(n231) );
  NAND2_X2 U358 ( .A1(\U7/DATA1_111 ), .A2(n1363), .ZN(n232) );
  NAND2_X2 U360 ( .A1(\U7/DATA1_110 ), .A2(n1363), .ZN(n233) );
  NAND2_X2 U362 ( .A1(\U7/DATA1_11 ), .A2(n1364), .ZN(n234) );
  NAND2_X2 U364 ( .A1(\U7/DATA1_109 ), .A2(n1363), .ZN(n235) );
  NAND2_X2 U366 ( .A1(\U7/DATA1_108 ), .A2(n1363), .ZN(n236) );
  NAND2_X2 U368 ( .A1(\U7/DATA1_107 ), .A2(n1363), .ZN(n237) );
  NAND2_X2 U370 ( .A1(\U7/DATA1_106 ), .A2(n1363), .ZN(n238) );
  NAND2_X2 U372 ( .A1(\U7/DATA1_105 ), .A2(n1363), .ZN(n239) );
  NAND2_X2 U374 ( .A1(\U7/DATA1_104 ), .A2(n1363), .ZN(n240) );
  NAND2_X2 U376 ( .A1(\U7/DATA1_103 ), .A2(n1363), .ZN(n241) );
  NAND2_X2 U378 ( .A1(\U7/DATA1_102 ), .A2(n1363), .ZN(n242) );
  NAND2_X2 U380 ( .A1(\U7/DATA1_101 ), .A2(n1363), .ZN(n243) );
  NAND2_X2 U382 ( .A1(\U7/DATA1_100 ), .A2(n1363), .ZN(n244) );
  NAND2_X2 U385 ( .A1(\U7/DATA1_10 ), .A2(n1364), .ZN(n245) );
  NAND2_X2 U387 ( .A1(\U7/DATA1_1 ), .A2(n1364), .ZN(n246) );
  NAND2_X2 U389 ( .A1(\U7/DATA1_0 ), .A2(n1364), .ZN(n247) );
  NAND2_X2 U391 ( .A1(PosElement[0]), .A2(PosElement[1]), .ZN(n62) );
  INV_X4 U3 ( .A(1'b0), .ZN(RowReady) );
  NAND2_X4 U7 ( .A1(PosElement[1]), .A2(n1436), .ZN(n1363) );
  NAND2_X4 U9 ( .A1(PosElement[1]), .A2(n50), .ZN(n1364) );
  OR2_X4 U11 ( .A1(n1485), .A2(PosElement[0]), .ZN(n50) );
  AND3_X4 U13 ( .A1(n50), .A2(n62), .A3(n1432), .ZN(n1365) );
  INV_X4 U15 ( .A(n1365), .ZN(n1434) );
  INV_X4 U17 ( .A(n1365), .ZN(n1433) );
  INV_X4 U19 ( .A(n1430), .ZN(n1432) );
  INV_X4 U21 ( .A(n1435), .ZN(n1436) );
  INV_X4 U23 ( .A(n1430), .ZN(n1431) );
  OAI21_X2 U25 ( .B1(n50), .B2(n1484), .A(n92), .ZN(\U4/Z_64 ) );
  OAI21_X2 U27 ( .B1(n50), .B2(n1483), .A(n91), .ZN(\U4/Z_65 ) );
  OAI21_X2 U29 ( .B1(n50), .B2(n1482), .A(n90), .ZN(\U4/Z_66 ) );
  OAI21_X2 U31 ( .B1(n50), .B2(n1481), .A(n89), .ZN(\U4/Z_67 ) );
  OAI21_X2 U33 ( .B1(n50), .B2(n1480), .A(n88), .ZN(\U4/Z_68 ) );
  OAI21_X2 U35 ( .B1(n50), .B2(n1479), .A(n87), .ZN(\U4/Z_69 ) );
  OAI21_X2 U37 ( .B1(n50), .B2(n1478), .A(n85), .ZN(\U4/Z_70 ) );
  OAI21_X2 U39 ( .B1(n50), .B2(n1477), .A(n84), .ZN(\U4/Z_71 ) );
  OAI21_X2 U41 ( .B1(n50), .B2(n1476), .A(n83), .ZN(\U4/Z_72 ) );
  OAI21_X2 U43 ( .B1(n50), .B2(n1475), .A(n82), .ZN(\U4/Z_73 ) );
  OAI21_X2 U45 ( .B1(n50), .B2(n1474), .A(n81), .ZN(\U4/Z_74 ) );
  OAI21_X2 U47 ( .B1(n50), .B2(n1468), .A(n74), .ZN(\U4/Z_80 ) );
  OAI21_X2 U49 ( .B1(n50), .B2(n1467), .A(n73), .ZN(\U4/Z_81 ) );
  OAI21_X2 U51 ( .B1(n50), .B2(n1466), .A(n72), .ZN(\U4/Z_82 ) );
  OAI21_X2 U53 ( .B1(n50), .B2(n1465), .A(n71), .ZN(\U4/Z_83 ) );
  OAI21_X2 U55 ( .B1(n50), .B2(n1464), .A(n70), .ZN(\U4/Z_84 ) );
  OAI21_X2 U57 ( .B1(n50), .B2(n1463), .A(n69), .ZN(\U4/Z_85 ) );
  OAI21_X2 U59 ( .B1(n50), .B2(n1462), .A(n68), .ZN(\U4/Z_86 ) );
  OAI21_X2 U61 ( .B1(n50), .B2(n1461), .A(n67), .ZN(\U4/Z_87 ) );
  OAI21_X2 U63 ( .B1(n50), .B2(n1460), .A(n66), .ZN(\U4/Z_88 ) );
  OAI21_X2 U65 ( .B1(n50), .B2(n1459), .A(n65), .ZN(\U4/Z_89 ) );
  OAI21_X2 U67 ( .B1(n50), .B2(n1448), .A(n244), .ZN(\U4/Z_100 ) );
  OAI21_X2 U69 ( .B1(n50), .B2(n1447), .A(n243), .ZN(\U4/Z_101 ) );
  OAI21_X2 U71 ( .B1(n50), .B2(n1446), .A(n242), .ZN(\U4/Z_102 ) );
  OAI21_X2 U73 ( .B1(n50), .B2(n1445), .A(n241), .ZN(\U4/Z_103 ) );
  OAI21_X2 U75 ( .B1(n50), .B2(n1444), .A(n240), .ZN(\U4/Z_104 ) );
  OAI21_X2 U77 ( .B1(n50), .B2(n1443), .A(n239), .ZN(\U4/Z_105 ) );
  OAI21_X2 U79 ( .B1(n50), .B2(n1442), .A(n238), .ZN(\U4/Z_106 ) );
  OAI21_X2 U81 ( .B1(n50), .B2(n1458), .A(n61), .ZN(\U4/Z_90 ) );
  OAI21_X2 U83 ( .B1(n50), .B2(n1452), .A(n55), .ZN(\U4/Z_96 ) );
  OAI21_X2 U85 ( .B1(n50), .B2(n1451), .A(n54), .ZN(\U4/Z_97 ) );
  OAI21_X2 U87 ( .B1(n50), .B2(n1450), .A(n53), .ZN(\U4/Z_98 ) );
  OAI21_X2 U89 ( .B1(n50), .B2(n1449), .A(n51), .ZN(\U4/Z_99 ) );
  INV_X4 U91 ( .A(n62), .ZN(n1435) );
  INV_X4 U93 ( .A(n175), .ZN(n1430) );
  BUF_X4 U95 ( .A(\U4/Z_48 ), .Z(PaddedRow[48]) );
  BUF_X4 U97 ( .A(\U4/Z_49 ), .Z(PaddedRow[49]) );
  BUF_X4 U99 ( .A(\U4/Z_50 ), .Z(PaddedRow[50]) );
  BUF_X4 U101 ( .A(\U4/Z_51 ), .Z(PaddedRow[51]) );
  BUF_X4 U103 ( .A(\U4/Z_52 ), .Z(PaddedRow[52]) );
  BUF_X4 U105 ( .A(\U4/Z_53 ), .Z(PaddedRow[53]) );
  BUF_X4 U107 ( .A(\U4/Z_54 ), .Z(PaddedRow[54]) );
  BUF_X4 U109 ( .A(\U4/Z_55 ), .Z(PaddedRow[55]) );
  BUF_X4 U111 ( .A(\U4/Z_56 ), .Z(PaddedRow[56]) );
  BUF_X4 U113 ( .A(\U4/Z_57 ), .Z(PaddedRow[57]) );
  BUF_X4 U115 ( .A(\U4/Z_58 ), .Z(PaddedRow[58]) );
  BUF_X4 U117 ( .A(\U4/Z_59 ), .Z(PaddedRow[59]) );
  BUF_X4 U119 ( .A(\U4/Z_60 ), .Z(PaddedRow[60]) );
  BUF_X4 U121 ( .A(\U4/Z_61 ), .Z(PaddedRow[61]) );
  BUF_X4 U123 ( .A(\U4/Z_62 ), .Z(PaddedRow[62]) );
  BUF_X4 U125 ( .A(\U4/Z_63 ), .Z(PaddedRow[63]) );
  BUF_X4 U127 ( .A(\U4/Z_112 ), .Z(PaddedRow[112]) );
  BUF_X4 U129 ( .A(\U4/Z_113 ), .Z(PaddedRow[113]) );
  BUF_X4 U131 ( .A(\U4/Z_114 ), .Z(PaddedRow[114]) );
  BUF_X4 U133 ( .A(\U4/Z_115 ), .Z(PaddedRow[115]) );
  BUF_X4 U135 ( .A(\U4/Z_116 ), .Z(PaddedRow[116]) );
  BUF_X4 U137 ( .A(\U4/Z_117 ), .Z(PaddedRow[117]) );
  BUF_X4 U139 ( .A(\U4/Z_118 ), .Z(PaddedRow[118]) );
  BUF_X4 U141 ( .A(\U4/Z_119 ), .Z(PaddedRow[119]) );
  BUF_X4 U143 ( .A(\U4/Z_120 ), .Z(PaddedRow[120]) );
  BUF_X4 U145 ( .A(\U4/Z_121 ), .Z(PaddedRow[121]) );
  BUF_X4 U147 ( .A(\U4/Z_122 ), .Z(PaddedRow[122]) );
  BUF_X4 U149 ( .A(\U4/Z_123 ), .Z(PaddedRow[123]) );
  BUF_X4 U151 ( .A(\U4/Z_124 ), .Z(PaddedRow[124]) );
  BUF_X4 U153 ( .A(\U4/Z_125 ), .Z(PaddedRow[125]) );
  BUF_X4 U155 ( .A(\U4/Z_126 ), .Z(PaddedRow[126]) );
  BUF_X4 U157 ( .A(\U4/Z_127 ), .Z(PaddedRow[127]) );
  BUF_X4 U159 ( .A(\U4/Z_176 ), .Z(PaddedRow[176]) );
  BUF_X4 U161 ( .A(\U4/Z_177 ), .Z(PaddedRow[177]) );
  BUF_X4 U163 ( .A(\U4/Z_178 ), .Z(PaddedRow[178]) );
  BUF_X4 U165 ( .A(\U4/Z_179 ), .Z(PaddedRow[179]) );
  BUF_X4 U167 ( .A(\U4/Z_180 ), .Z(PaddedRow[180]) );
  BUF_X4 U169 ( .A(\U4/Z_181 ), .Z(PaddedRow[181]) );
  BUF_X4 U171 ( .A(\U4/Z_182 ), .Z(PaddedRow[182]) );
  BUF_X4 U173 ( .A(\U4/Z_183 ), .Z(PaddedRow[183]) );
  BUF_X4 U175 ( .A(\U4/Z_184 ), .Z(PaddedRow[184]) );
  BUF_X4 U177 ( .A(\U4/Z_185 ), .Z(PaddedRow[185]) );
  BUF_X4 U179 ( .A(\U4/Z_186 ), .Z(PaddedRow[186]) );
  BUF_X4 U181 ( .A(\U4/Z_187 ), .Z(PaddedRow[187]) );
  BUF_X4 U183 ( .A(\U4/Z_188 ), .Z(PaddedRow[188]) );
  BUF_X4 U185 ( .A(\U4/Z_189 ), .Z(PaddedRow[189]) );
  BUF_X4 U187 ( .A(\U4/Z_190 ), .Z(PaddedRow[190]) );
  BUF_X4 U189 ( .A(\U4/Z_191 ), .Z(PaddedRow[191]) );
  BUF_X4 U191 ( .A(\U4/Z_240 ), .Z(PaddedRow[240]) );
  BUF_X4 U193 ( .A(\U4/Z_241 ), .Z(PaddedRow[241]) );
  BUF_X4 U195 ( .A(\U4/Z_242 ), .Z(PaddedRow[242]) );
  BUF_X4 U197 ( .A(\U4/Z_243 ), .Z(PaddedRow[243]) );
  BUF_X4 U199 ( .A(\U4/Z_244 ), .Z(PaddedRow[244]) );
  BUF_X4 U201 ( .A(\U4/Z_245 ), .Z(PaddedRow[245]) );
  BUF_X4 U203 ( .A(\U4/Z_246 ), .Z(PaddedRow[246]) );
  BUF_X4 U205 ( .A(\U4/Z_247 ), .Z(PaddedRow[247]) );
  BUF_X4 U207 ( .A(\U4/Z_248 ), .Z(PaddedRow[248]) );
  BUF_X4 U209 ( .A(\U4/Z_249 ), .Z(PaddedRow[249]) );
  BUF_X4 U211 ( .A(\U4/Z_250 ), .Z(PaddedRow[250]) );
  BUF_X4 U213 ( .A(\U4/Z_251 ), .Z(PaddedRow[251]) );
  BUF_X4 U215 ( .A(\U4/Z_252 ), .Z(PaddedRow[252]) );
  BUF_X4 U217 ( .A(\U4/Z_253 ), .Z(PaddedRow[253]) );
  BUF_X4 U219 ( .A(\U4/Z_254 ), .Z(PaddedRow[254]) );
  BUF_X4 U221 ( .A(\U4/Z_255 ), .Z(PaddedRow[255]) );
  OAI21_X2 U223 ( .B1(n1436), .B2(n1484), .A(n247), .ZN(\U4/Z_0 ) );
  OAI21_X2 U225 ( .B1(n1436), .B2(n1483), .A(n246), .ZN(\U4/Z_1 ) );
  OAI21_X2 U227 ( .B1(n1436), .B2(n1482), .A(n166), .ZN(\U4/Z_2 ) );
  OAI21_X2 U229 ( .B1(n1436), .B2(n1481), .A(n114), .ZN(\U4/Z_3 ) );
  OAI21_X2 U231 ( .B1(n1436), .B2(n1480), .A(n103), .ZN(\U4/Z_4 ) );
  OAI21_X2 U233 ( .B1(n1436), .B2(n1479), .A(n94), .ZN(\U4/Z_5 ) );
  OAI21_X2 U235 ( .B1(n1436), .B2(n1478), .A(n93), .ZN(\U4/Z_6 ) );
  OAI21_X2 U237 ( .B1(n1436), .B2(n1477), .A(n86), .ZN(\U4/Z_7 ) );
  OAI21_X2 U239 ( .B1(n1436), .B2(n1476), .A(n75), .ZN(\U4/Z_8 ) );
  OAI21_X2 U241 ( .B1(n62), .B2(n1475), .A(n63), .ZN(\U4/Z_9 ) );
  OAI21_X2 U243 ( .B1(n62), .B2(n1474), .A(n245), .ZN(\U4/Z_10 ) );
  OAI21_X2 U244 ( .B1(n62), .B2(n1473), .A(n234), .ZN(\U4/Z_11 ) );
  OAI21_X2 U246 ( .B1(n1436), .B2(n1472), .A(n231), .ZN(\U4/Z_12 ) );
  OAI21_X2 U248 ( .B1(n1436), .B2(n1471), .A(n228), .ZN(\U4/Z_13 ) );
  OAI21_X2 U250 ( .B1(n1436), .B2(n1470), .A(n217), .ZN(\U4/Z_14 ) );
  OAI21_X2 U252 ( .B1(n1436), .B2(n1469), .A(n206), .ZN(\U4/Z_15 ) );
  OAI21_X2 U254 ( .B1(n1436), .B2(n1468), .A(n195), .ZN(\U4/Z_16 ) );
  OAI21_X2 U256 ( .B1(n1436), .B2(n1467), .A(n184), .ZN(\U4/Z_17 ) );
  OAI21_X2 U258 ( .B1(n1436), .B2(n1466), .A(n177), .ZN(\U4/Z_18 ) );
  OAI21_X2 U260 ( .B1(n1436), .B2(n1465), .A(n176), .ZN(\U4/Z_19 ) );
  OAI21_X2 U262 ( .B1(n1436), .B2(n1464), .A(n165), .ZN(\U4/Z_20 ) );
  OAI21_X2 U264 ( .B1(n62), .B2(n1463), .A(n154), .ZN(\U4/Z_21 ) );
  OAI21_X2 U266 ( .B1(n1436), .B2(n1462), .A(n143), .ZN(\U4/Z_22 ) );
  OAI21_X2 U268 ( .B1(n1436), .B2(n1461), .A(n132), .ZN(\U4/Z_23 ) );
  OAI21_X2 U270 ( .B1(n62), .B2(n1460), .A(n120), .ZN(\U4/Z_24 ) );
  OAI21_X2 U272 ( .B1(n62), .B2(n1459), .A(n119), .ZN(\U4/Z_25 ) );
  OAI21_X2 U274 ( .B1(n1458), .B2(n1436), .A(n118), .ZN(\U4/Z_26 ) );
  OAI21_X2 U276 ( .B1(n1457), .B2(n62), .A(n117), .ZN(\U4/Z_27 ) );
  OAI21_X2 U278 ( .B1(n1456), .B2(n62), .A(n116), .ZN(\U4/Z_28 ) );
  OAI21_X2 U280 ( .B1(n1455), .B2(n62), .A(n115), .ZN(\U4/Z_29 ) );
  OAI21_X2 U282 ( .B1(n1454), .B2(n62), .A(n113), .ZN(\U4/Z_30 ) );
  OAI21_X2 U284 ( .B1(n1453), .B2(n62), .A(n112), .ZN(\U4/Z_31 ) );
  OAI21_X2 U286 ( .B1(n1452), .B2(n62), .A(n111), .ZN(\U4/Z_32 ) );
  OAI21_X2 U288 ( .B1(n1451), .B2(n62), .A(n110), .ZN(\U4/Z_33 ) );
  OAI21_X2 U290 ( .B1(n1450), .B2(n62), .A(n109), .ZN(\U4/Z_34 ) );
  OAI21_X2 U292 ( .B1(n1449), .B2(n62), .A(n108), .ZN(\U4/Z_35 ) );
  OAI21_X2 U294 ( .B1(n62), .B2(n1448), .A(n107), .ZN(\U4/Z_36 ) );
  OAI21_X2 U296 ( .B1(n62), .B2(n1447), .A(n106), .ZN(\U4/Z_37 ) );
  OAI21_X2 U298 ( .B1(n62), .B2(n1446), .A(n105), .ZN(\U4/Z_38 ) );
  OAI21_X2 U300 ( .B1(n62), .B2(n1445), .A(n104), .ZN(\U4/Z_39 ) );
  OAI21_X2 U302 ( .B1(n62), .B2(n1444), .A(n102), .ZN(\U4/Z_40 ) );
  OAI21_X2 U304 ( .B1(n1436), .B2(n1443), .A(n101), .ZN(\U4/Z_41 ) );
  OAI21_X2 U306 ( .B1(n1436), .B2(n1442), .A(n100), .ZN(\U4/Z_42 ) );
  OAI21_X2 U308 ( .B1(n1436), .B2(n1441), .A(n99), .ZN(\U4/Z_43 ) );
  OAI21_X2 U310 ( .B1(n1436), .B2(n1440), .A(n98), .ZN(\U4/Z_44 ) );
  OAI21_X2 U312 ( .B1(n1436), .B2(n1439), .A(n97), .ZN(\U4/Z_45 ) );
  OAI21_X2 U314 ( .B1(n1436), .B2(n1438), .A(n96), .ZN(\U4/Z_46 ) );
  OAI21_X2 U316 ( .B1(n1436), .B2(n1437), .A(n95), .ZN(\U4/Z_47 ) );
  OAI21_X2 U318 ( .B1(n50), .B2(n1473), .A(n80), .ZN(\U4/Z_75 ) );
  OAI21_X2 U320 ( .B1(n50), .B2(n1472), .A(n79), .ZN(\U4/Z_76 ) );
  OAI21_X2 U322 ( .B1(n50), .B2(n1471), .A(n78), .ZN(\U4/Z_77 ) );
  OAI21_X2 U324 ( .B1(n50), .B2(n1470), .A(n77), .ZN(\U4/Z_78 ) );
  OAI21_X2 U326 ( .B1(n50), .B2(n1469), .A(n76), .ZN(\U4/Z_79 ) );
  OAI21_X2 U328 ( .B1(n50), .B2(n1441), .A(n237), .ZN(\U4/Z_107 ) );
  OAI21_X2 U330 ( .B1(n50), .B2(n1440), .A(n236), .ZN(\U4/Z_108 ) );
  OAI21_X2 U332 ( .B1(n50), .B2(n1439), .A(n235), .ZN(\U4/Z_109 ) );
  OAI21_X2 U334 ( .B1(n50), .B2(n1438), .A(n233), .ZN(\U4/Z_110 ) );
  OAI21_X2 U336 ( .B1(n50), .B2(n1437), .A(n232), .ZN(\U4/Z_111 ) );
  OAI21_X2 U338 ( .B1(n1484), .B2(n1433), .A(n174), .ZN(\U4/Z_192 ) );
  OAI21_X2 U340 ( .B1(n1483), .B2(n1433), .A(n173), .ZN(\U4/Z_193 ) );
  OAI21_X2 U342 ( .B1(n1482), .B2(n1433), .A(n172), .ZN(\U4/Z_194 ) );
  OAI21_X2 U344 ( .B1(n1481), .B2(n1433), .A(n171), .ZN(\U4/Z_195 ) );
  OAI21_X2 U346 ( .B1(n1480), .B2(n1433), .A(n170), .ZN(\U4/Z_196 ) );
  OAI21_X2 U348 ( .B1(n1479), .B2(n1433), .A(n169), .ZN(\U4/Z_197 ) );
  OAI21_X2 U350 ( .B1(n1478), .B2(n1433), .A(n168), .ZN(\U4/Z_198 ) );
  OAI21_X2 U352 ( .B1(n1477), .B2(n1433), .A(n167), .ZN(\U4/Z_199 ) );
  OAI21_X2 U355 ( .B1(n1476), .B2(n1433), .A(n164), .ZN(\U4/Z_200 ) );
  OAI21_X2 U357 ( .B1(n1475), .B2(n1433), .A(n163), .ZN(\U4/Z_201 ) );
  OAI21_X2 U359 ( .B1(n1474), .B2(n1433), .A(n162), .ZN(\U4/Z_202 ) );
  OAI21_X2 U361 ( .B1(n1473), .B2(n1433), .A(n161), .ZN(\U4/Z_203 ) );
  OAI21_X2 U363 ( .B1(n1472), .B2(n1434), .A(n160), .ZN(\U4/Z_204 ) );
  OAI21_X2 U365 ( .B1(n1471), .B2(n1433), .A(n159), .ZN(\U4/Z_205 ) );
  OAI21_X2 U367 ( .B1(n1470), .B2(n1433), .A(n158), .ZN(\U4/Z_206 ) );
  OAI21_X2 U369 ( .B1(n1469), .B2(n1433), .A(n157), .ZN(\U4/Z_207 ) );
  OAI21_X2 U371 ( .B1(n1468), .B2(n1433), .A(n156), .ZN(\U4/Z_208 ) );
  OAI21_X2 U373 ( .B1(n1467), .B2(n1433), .A(n155), .ZN(\U4/Z_209 ) );
  OAI21_X2 U375 ( .B1(n1466), .B2(n1434), .A(n153), .ZN(\U4/Z_210 ) );
  OAI21_X2 U377 ( .B1(n1465), .B2(n1433), .A(n152), .ZN(\U4/Z_211 ) );
  OAI21_X2 U379 ( .B1(n1464), .B2(n1433), .A(n151), .ZN(\U4/Z_212 ) );
  OAI21_X2 U381 ( .B1(n1463), .B2(n1434), .A(n150), .ZN(\U4/Z_213 ) );
  OAI21_X2 U383 ( .B1(n1462), .B2(n1433), .A(n149), .ZN(\U4/Z_214 ) );
  OAI21_X2 U384 ( .B1(n1461), .B2(n1433), .A(n148), .ZN(\U4/Z_215 ) );
  OAI21_X2 U386 ( .B1(n1460), .B2(n1433), .A(n147), .ZN(\U4/Z_216 ) );
  OAI21_X2 U388 ( .B1(n1459), .B2(n1434), .A(n146), .ZN(\U4/Z_217 ) );
  OAI21_X2 U390 ( .B1(n1458), .B2(n1433), .A(n145), .ZN(\U4/Z_218 ) );
  OAI21_X2 U392 ( .B1(n1457), .B2(n1433), .A(n144), .ZN(\U4/Z_219 ) );
  OAI21_X2 U393 ( .B1(n1456), .B2(n1433), .A(n142), .ZN(\U4/Z_220 ) );
  OAI21_X2 U394 ( .B1(n1455), .B2(n1433), .A(n141), .ZN(\U4/Z_221 ) );
  OAI21_X2 U395 ( .B1(n1454), .B2(n1433), .A(n140), .ZN(\U4/Z_222 ) );
  OAI21_X2 U396 ( .B1(n1453), .B2(n1433), .A(n139), .ZN(\U4/Z_223 ) );
  OAI21_X2 U397 ( .B1(n1452), .B2(n1433), .A(n138), .ZN(\U4/Z_224 ) );
  OAI21_X2 U398 ( .B1(n1451), .B2(n1433), .A(n137), .ZN(\U4/Z_225 ) );
  OAI21_X2 U399 ( .B1(n1450), .B2(n1433), .A(n136), .ZN(\U4/Z_226 ) );
  OAI21_X2 U400 ( .B1(n1449), .B2(n1433), .A(n135), .ZN(\U4/Z_227 ) );
  OAI21_X2 U401 ( .B1(n1448), .B2(n1433), .A(n134), .ZN(\U4/Z_228 ) );
  OAI21_X2 U402 ( .B1(n1447), .B2(n1433), .A(n133), .ZN(\U4/Z_229 ) );
  OAI21_X2 U403 ( .B1(n1446), .B2(n1433), .A(n131), .ZN(\U4/Z_230 ) );
  OAI21_X2 U404 ( .B1(n1445), .B2(n1433), .A(n130), .ZN(\U4/Z_231 ) );
  OAI21_X2 U405 ( .B1(n1444), .B2(n1433), .A(n129), .ZN(\U4/Z_232 ) );
  OAI21_X2 U406 ( .B1(n1443), .B2(n1433), .A(n128), .ZN(\U4/Z_233 ) );
  OAI21_X2 U407 ( .B1(n1442), .B2(n1433), .A(n127), .ZN(\U4/Z_234 ) );
  OAI21_X2 U408 ( .B1(n1441), .B2(n1434), .A(n126), .ZN(\U4/Z_235 ) );
  OAI21_X2 U409 ( .B1(n1440), .B2(n1433), .A(n125), .ZN(\U4/Z_236 ) );
  OAI21_X2 U410 ( .B1(n1439), .B2(n1433), .A(n124), .ZN(\U4/Z_237 ) );
  OAI21_X2 U411 ( .B1(n1438), .B2(n1433), .A(n123), .ZN(\U4/Z_238 ) );
  OAI21_X2 U412 ( .B1(n1437), .B2(n1434), .A(n122), .ZN(\U4/Z_239 ) );
  OAI21_X2 U413 ( .B1(n50), .B2(n1457), .A(n60), .ZN(\U4/Z_91 ) );
  OAI21_X2 U414 ( .B1(n50), .B2(n1456), .A(n59), .ZN(\U4/Z_92 ) );
  OAI21_X2 U415 ( .B1(n50), .B2(n1455), .A(n58), .ZN(\U4/Z_93 ) );
  OAI21_X2 U416 ( .B1(n50), .B2(n1454), .A(n57), .ZN(\U4/Z_94 ) );
  OAI21_X2 U417 ( .B1(n50), .B2(n1453), .A(n56), .ZN(\U4/Z_95 ) );
  OAI21_X2 U418 ( .B1(n1484), .B2(n1431), .A(n230), .ZN(\U4/Z_128 ) );
  OAI21_X2 U419 ( .B1(n1483), .B2(n1431), .A(n229), .ZN(\U4/Z_129 ) );
  OAI21_X2 U420 ( .B1(n1482), .B2(n1431), .A(n227), .ZN(\U4/Z_130 ) );
  OAI21_X2 U421 ( .B1(n1481), .B2(n1431), .A(n226), .ZN(\U4/Z_131 ) );
  OAI21_X2 U422 ( .B1(n1480), .B2(n1431), .A(n225), .ZN(\U4/Z_132 ) );
  OAI21_X2 U423 ( .B1(n1479), .B2(n1431), .A(n224), .ZN(\U4/Z_133 ) );
  OAI21_X2 U424 ( .B1(n1478), .B2(n1431), .A(n223), .ZN(\U4/Z_134 ) );
  OAI21_X2 U425 ( .B1(n1477), .B2(n1431), .A(n222), .ZN(\U4/Z_135 ) );
  OAI21_X2 U426 ( .B1(n1476), .B2(n1431), .A(n221), .ZN(\U4/Z_136 ) );
  OAI21_X2 U427 ( .B1(n1475), .B2(n1431), .A(n220), .ZN(\U4/Z_137 ) );
  OAI21_X2 U428 ( .B1(n1474), .B2(n1431), .A(n219), .ZN(\U4/Z_138 ) );
  OAI21_X2 U429 ( .B1(n1473), .B2(n1431), .A(n218), .ZN(\U4/Z_139 ) );
  OAI21_X2 U430 ( .B1(n1472), .B2(n1431), .A(n216), .ZN(\U4/Z_140 ) );
  OAI21_X2 U431 ( .B1(n1471), .B2(n1431), .A(n215), .ZN(\U4/Z_141 ) );
  OAI21_X2 U432 ( .B1(n1470), .B2(n1431), .A(n214), .ZN(\U4/Z_142 ) );
  OAI21_X2 U433 ( .B1(n1469), .B2(n1431), .A(n213), .ZN(\U4/Z_143 ) );
  OAI21_X2 U434 ( .B1(n1468), .B2(n1431), .A(n212), .ZN(\U4/Z_144 ) );
  OAI21_X2 U435 ( .B1(n1467), .B2(n1431), .A(n211), .ZN(\U4/Z_145 ) );
  OAI21_X2 U436 ( .B1(n1466), .B2(n1431), .A(n210), .ZN(\U4/Z_146 ) );
  OAI21_X2 U437 ( .B1(n1465), .B2(n1431), .A(n209), .ZN(\U4/Z_147 ) );
  OAI21_X2 U438 ( .B1(n1464), .B2(n1431), .A(n208), .ZN(\U4/Z_148 ) );
  OAI21_X2 U439 ( .B1(n1463), .B2(n1431), .A(n207), .ZN(\U4/Z_149 ) );
  OAI21_X2 U440 ( .B1(n1462), .B2(n1431), .A(n205), .ZN(\U4/Z_150 ) );
  OAI21_X2 U441 ( .B1(n1461), .B2(n1431), .A(n204), .ZN(\U4/Z_151 ) );
  OAI21_X2 U442 ( .B1(n1460), .B2(n1431), .A(n203), .ZN(\U4/Z_152 ) );
  OAI21_X2 U443 ( .B1(n1459), .B2(n1431), .A(n202), .ZN(\U4/Z_153 ) );
  OAI21_X2 U444 ( .B1(n1458), .B2(n1431), .A(n201), .ZN(\U4/Z_154 ) );
  OAI21_X2 U445 ( .B1(n1457), .B2(n1431), .A(n200), .ZN(\U4/Z_155 ) );
  OAI21_X2 U446 ( .B1(n1456), .B2(n1431), .A(n199), .ZN(\U4/Z_156 ) );
  OAI21_X2 U447 ( .B1(n1455), .B2(n1431), .A(n198), .ZN(\U4/Z_157 ) );
  OAI21_X2 U448 ( .B1(n1454), .B2(n1431), .A(n197), .ZN(\U4/Z_158 ) );
  OAI21_X2 U449 ( .B1(n1453), .B2(n1431), .A(n196), .ZN(\U4/Z_159 ) );
  OAI21_X2 U450 ( .B1(n1452), .B2(n1431), .A(n194), .ZN(\U4/Z_160 ) );
  OAI21_X2 U451 ( .B1(n1451), .B2(n1431), .A(n193), .ZN(\U4/Z_161 ) );
  OAI21_X2 U452 ( .B1(n1450), .B2(n1431), .A(n192), .ZN(\U4/Z_162 ) );
  OAI21_X2 U453 ( .B1(n1449), .B2(n1431), .A(n191), .ZN(\U4/Z_163 ) );
  OAI21_X2 U454 ( .B1(n1448), .B2(n1431), .A(n190), .ZN(\U4/Z_164 ) );
  OAI21_X2 U455 ( .B1(n1447), .B2(n1431), .A(n189), .ZN(\U4/Z_165 ) );
  OAI21_X2 U456 ( .B1(n1446), .B2(n1431), .A(n188), .ZN(\U4/Z_166 ) );
  OAI21_X2 U457 ( .B1(n1445), .B2(n1431), .A(n187), .ZN(\U4/Z_167 ) );
  OAI21_X2 U458 ( .B1(n1444), .B2(n1431), .A(n186), .ZN(\U4/Z_168 ) );
  OAI21_X2 U459 ( .B1(n1443), .B2(n1431), .A(n185), .ZN(\U4/Z_169 ) );
  OAI21_X2 U460 ( .B1(n1442), .B2(n1431), .A(n183), .ZN(\U4/Z_170 ) );
  OAI21_X2 U461 ( .B1(n1441), .B2(n1431), .A(n182), .ZN(\U4/Z_171 ) );
  OAI21_X2 U462 ( .B1(n1440), .B2(n1431), .A(n181), .ZN(\U4/Z_172 ) );
  OAI21_X2 U463 ( .B1(n1439), .B2(n1431), .A(n180), .ZN(\U4/Z_173 ) );
  OAI21_X2 U464 ( .B1(n1438), .B2(n1431), .A(n179), .ZN(\U4/Z_174 ) );
  OAI21_X2 U465 ( .B1(n1437), .B2(n1431), .A(n178), .ZN(\U4/Z_175 ) );
  INV_X4 U466 ( .A(\U7/DATA1_239 ), .ZN(n1437) );
  INV_X4 U467 ( .A(\U7/DATA1_238 ), .ZN(n1438) );
  INV_X4 U468 ( .A(\U7/DATA1_237 ), .ZN(n1439) );
  INV_X4 U469 ( .A(\U7/DATA1_236 ), .ZN(n1440) );
  INV_X4 U470 ( .A(\U7/DATA1_235 ), .ZN(n1441) );
  INV_X4 U471 ( .A(\U7/DATA1_234 ), .ZN(n1442) );
  INV_X4 U472 ( .A(\U7/DATA1_233 ), .ZN(n1443) );
  INV_X4 U473 ( .A(\U7/DATA1_232 ), .ZN(n1444) );
  INV_X4 U474 ( .A(\U7/DATA1_231 ), .ZN(n1445) );
  INV_X4 U475 ( .A(\U7/DATA1_230 ), .ZN(n1446) );
  INV_X4 U476 ( .A(\U7/DATA1_229 ), .ZN(n1447) );
  INV_X4 U477 ( .A(\U7/DATA1_228 ), .ZN(n1448) );
  INV_X4 U478 ( .A(\U7/DATA1_227 ), .ZN(n1449) );
  INV_X4 U479 ( .A(\U7/DATA1_226 ), .ZN(n1450) );
  INV_X4 U480 ( .A(\U7/DATA1_225 ), .ZN(n1451) );
  INV_X4 U481 ( .A(\U7/DATA1_224 ), .ZN(n1452) );
  INV_X4 U482 ( .A(\U7/DATA1_223 ), .ZN(n1453) );
  INV_X4 U483 ( .A(\U7/DATA1_222 ), .ZN(n1454) );
  INV_X4 U484 ( .A(\U7/DATA1_221 ), .ZN(n1455) );
  INV_X4 U485 ( .A(\U7/DATA1_220 ), .ZN(n1456) );
  INV_X4 U486 ( .A(\U7/DATA1_219 ), .ZN(n1457) );
  INV_X4 U487 ( .A(\U7/DATA1_218 ), .ZN(n1458) );
  INV_X4 U488 ( .A(\U7/DATA1_217 ), .ZN(n1459) );
  INV_X4 U489 ( .A(\U7/DATA1_216 ), .ZN(n1460) );
  INV_X4 U490 ( .A(\U7/DATA1_215 ), .ZN(n1461) );
  INV_X4 U491 ( .A(\U7/DATA1_214 ), .ZN(n1462) );
  INV_X4 U492 ( .A(\U7/DATA1_213 ), .ZN(n1463) );
  INV_X4 U493 ( .A(\U7/DATA1_212 ), .ZN(n1464) );
  INV_X4 U494 ( .A(\U7/DATA1_211 ), .ZN(n1465) );
  INV_X4 U495 ( .A(\U7/DATA1_210 ), .ZN(n1466) );
  INV_X4 U496 ( .A(\U7/DATA1_209 ), .ZN(n1467) );
  INV_X4 U497 ( .A(\U7/DATA1_208 ), .ZN(n1468) );
  INV_X4 U498 ( .A(\U7/DATA1_207 ), .ZN(n1469) );
  INV_X4 U499 ( .A(\U7/DATA1_206 ), .ZN(n1470) );
  INV_X4 U500 ( .A(\U7/DATA1_205 ), .ZN(n1471) );
  INV_X4 U501 ( .A(\U7/DATA1_204 ), .ZN(n1472) );
  INV_X4 U502 ( .A(\U7/DATA1_203 ), .ZN(n1473) );
  INV_X4 U503 ( .A(\U7/DATA1_202 ), .ZN(n1474) );
  INV_X4 U504 ( .A(\U7/DATA1_201 ), .ZN(n1475) );
  INV_X4 U505 ( .A(\U7/DATA1_200 ), .ZN(n1476) );
  INV_X4 U506 ( .A(\U7/DATA1_199 ), .ZN(n1477) );
  INV_X4 U507 ( .A(\U7/DATA1_198 ), .ZN(n1478) );
  INV_X4 U508 ( .A(\U7/DATA1_197 ), .ZN(n1479) );
  INV_X4 U509 ( .A(\U7/DATA1_196 ), .ZN(n1480) );
  INV_X4 U510 ( .A(\U7/DATA1_195 ), .ZN(n1481) );
  INV_X4 U511 ( .A(\U7/DATA1_194 ), .ZN(n1482) );
  INV_X4 U512 ( .A(\U7/DATA1_193 ), .ZN(n1483) );
  INV_X4 U513 ( .A(\U7/DATA1_192 ), .ZN(n1484) );
  INV_X4 U514 ( .A(PosElement[1]), .ZN(n1485) );
endmodule


module selector ( dataY, count, found1, found2, found3, found4, EOF );
  input [255:0] dataY;
  output [2:0] count;
  output found1, found2, found3, found4, EOF;
  wire   \U4/Z_0 , n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24;
  assign EOF = \U4/Z_0 ;

  INV_X4 U3 ( .A(n8), .ZN(found4) );
  INV_X4 U7 ( .A(n13), .ZN(found2) );
  NAND3_X2 U8 ( .A1(found3), .A2(n8), .A3(found1), .ZN(n12) );
  INV_X4 U9 ( .A(n10), .ZN(found1) );
  INV_X4 U10 ( .A(n14), .ZN(found3) );
  NAND2_X2 U11 ( .A1(n14), .A2(n10), .ZN(n11) );
  NAND2_X2 U12 ( .A1(n15), .A2(n16), .ZN(\U4/Z_0 ) );
  NOR3_X2 U14 ( .A1(dataY[122]), .A2(dataY[124]), .A3(dataY[123]), .ZN(n20) );
  NOR3_X2 U15 ( .A1(n14), .A2(dataY[121]), .A3(dataY[120]), .ZN(n19) );
  NAND3_X2 U16 ( .A1(dataY[126]), .A2(dataY[125]), .A3(dataY[127]), .ZN(n14)
         );
  NOR3_X2 U17 ( .A1(dataY[58]), .A2(dataY[60]), .A3(dataY[59]), .ZN(n18) );
  NOR3_X2 U18 ( .A1(n8), .A2(dataY[57]), .A3(dataY[56]), .ZN(n17) );
  NAND3_X2 U19 ( .A1(dataY[62]), .A2(dataY[61]), .A3(dataY[63]), .ZN(n8) );
  NOR3_X2 U21 ( .A1(dataY[250]), .A2(dataY[252]), .A3(dataY[251]), .ZN(n24) );
  NOR3_X2 U22 ( .A1(n10), .A2(dataY[249]), .A3(dataY[248]), .ZN(n23) );
  NAND3_X2 U23 ( .A1(dataY[254]), .A2(dataY[253]), .A3(dataY[255]), .ZN(n10)
         );
  NOR3_X2 U24 ( .A1(dataY[186]), .A2(dataY[188]), .A3(dataY[187]), .ZN(n22) );
  NOR3_X2 U25 ( .A1(n13), .A2(dataY[185]), .A3(dataY[184]), .ZN(n21) );
  NAND3_X2 U26 ( .A1(dataY[190]), .A2(dataY[189]), .A3(dataY[191]), .ZN(n13)
         );
  INV_X4 U4 ( .A(1'b1), .ZN(count[2]) );
  OAI21_X2 U6 ( .B1(found2), .B2(found3), .A(n9), .ZN(count[1]) );
  OAI21_X2 U13 ( .B1(found2), .B2(n8), .A(n10), .ZN(n9) );
  AOI21_X2 U20 ( .B1(n11), .B2(n12), .A(found2), .ZN(count[0]) );
  AOI22_X2 U27 ( .A1(n21), .A2(n22), .B1(n23), .B2(n24), .ZN(n15) );
  AOI22_X2 U28 ( .A1(n17), .A2(n18), .B1(n19), .B2(n20), .ZN(n16) );
endmodule


module EOF_reg ( clock, reset, EOF, OP, sig );
  input clock, reset, EOF;
  output OP, sig;
  wire   n44, \U4/DATA2_1 , \U4/DATA2_2 , \U4/DATA2_3 , \U4/DATA2_4 ,
         \add_24/carry[5] , \add_24/carry[4] , \add_24/carry[3] ,
         \add_24/carry[2] , \add_24/A[0] , \add_24/A[1] , \add_24/A[2] ,
         \add_24/A[3] , \add_24/A[4] , \add_24/A[5] , n3, n5, n7, n8, n9, n10,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n61, n62, n63, n64,
         n65;

  HA_X1 \add_24/U1_1_1  ( .A(\add_24/A[1] ), .B(\add_24/A[0] ), .CO(
        \add_24/carry[2] ), .S(\U4/DATA2_1 ) );
  HA_X1 \add_24/U1_1_2  ( .A(\add_24/A[2] ), .B(\add_24/carry[2] ), .CO(
        \add_24/carry[3] ), .S(\U4/DATA2_2 ) );
  HA_X1 \add_24/U1_1_3  ( .A(\add_24/A[3] ), .B(\add_24/carry[3] ), .CO(
        \add_24/carry[4] ), .S(\U4/DATA2_3 ) );
  HA_X1 \add_24/U1_1_4  ( .A(\add_24/A[4] ), .B(\add_24/carry[4] ), .CO(
        \add_24/carry[5] ), .S(\U4/DATA2_4 ) );
  DFF_X1 OPCheck_reg ( .D(n35), .CK(clock), .Q(n44) );
  DFF_X1 \count_reg[0]  ( .D(n33), .CK(clock), .Q(\add_24/A[0] ), .QN(n10) );
  DFF_X1 \count_reg[5]  ( .D(n34), .CK(clock), .Q(\add_24/A[5] ), .QN(n3) );
  DFF_X1 \count_reg[4]  ( .D(n29), .CK(clock), .Q(\add_24/A[4] ), .QN(n5) );
  DFF_X1 \count_reg[3]  ( .D(n30), .CK(clock), .Q(\add_24/A[3] ), .QN(n7) );
  DFF_X1 \count_reg[1]  ( .D(n32), .CK(clock), .Q(\add_24/A[1] ), .QN(n9) );
  NAND2_X2 U3 ( .A1(n12), .A2(n13), .ZN(n28) );
  NAND3_X2 U4 ( .A1(n61), .A2(n14), .A3(sig), .ZN(n12) );
  NAND4_X2 U5 ( .A1(n64), .A2(n10), .A3(n15), .A4(n9), .ZN(n14) );
  NOR2_X2 U6 ( .A1(\add_24/A[5] ), .A2(\add_24/A[3] ), .ZN(n15) );
  NAND2_X2 U8 ( .A1(\U4/DATA2_4 ), .A2(n62), .ZN(n18) );
  NAND2_X2 U10 ( .A1(\U4/DATA2_3 ), .A2(n62), .ZN(n19) );
  NAND2_X2 U12 ( .A1(\U4/DATA2_2 ), .A2(n62), .ZN(n20) );
  NAND2_X2 U14 ( .A1(\U4/DATA2_1 ), .A2(n62), .ZN(n21) );
  OAI22_X2 U15 ( .A1(n17), .A2(n10), .B1(\add_24/A[0] ), .B2(n22), .ZN(n33) );
  NAND3_X2 U17 ( .A1(n62), .A2(n3), .A3(\add_24/carry[5] ), .ZN(n24) );
  NAND3_X2 U19 ( .A1(n13), .A2(n65), .A3(n22), .ZN(n17) );
  OAI22_X2 U21 ( .A1(\add_24/A[4] ), .A2(\add_24/A[3] ), .B1(\add_24/A[1] ), 
        .B2(n16), .ZN(n25) );
  AND3_X2 U22 ( .A1(n44), .A2(n65), .A3(n13), .ZN(n26) );
  NAND4_X2 U23 ( .A1(\add_24/A[5] ), .A2(\add_24/A[3] ), .A3(n44), .A4(n27), 
        .ZN(n13) );
  NOR4_X2 U24 ( .A1(reset), .A2(\add_24/A[0] ), .A3(n16), .A4(n9), .ZN(n27) );
  NAND2_X2 U25 ( .A1(n8), .A2(n5), .ZN(n16) );
  OR2_X1 U31 ( .A1(n26), .A2(EOF), .ZN(n35) );
  DFF_X2 OP_reg ( .D(n28), .CK(clock), .Q(sig) );
  DFF_X2 \count_reg[2]  ( .D(n31), .CK(clock), .Q(\add_24/A[2] ), .QN(n8) );
  BUF_X4 U7 ( .A(sig), .Z(OP) );
  OAI211_X2 U9 ( .C1(n3), .C2(n25), .A(n65), .B(n44), .ZN(n22) );
  OAI21_X2 U11 ( .B1(n17), .B2(n8), .A(n20), .ZN(n31) );
  OAI21_X2 U13 ( .B1(n9), .B2(n17), .A(n21), .ZN(n32) );
  OAI21_X2 U16 ( .B1(n7), .B2(n17), .A(n19), .ZN(n30) );
  OAI21_X2 U18 ( .B1(n17), .B2(n5), .A(n18), .ZN(n29) );
  OAI21_X2 U20 ( .B1(n23), .B2(n3), .A(n24), .ZN(n34) );
  AOI21_X2 U26 ( .B1(n62), .B2(n63), .A(n61), .ZN(n23) );
  INV_X4 U27 ( .A(n17), .ZN(n61) );
  INV_X4 U28 ( .A(n22), .ZN(n62) );
  INV_X4 U29 ( .A(\add_24/carry[5] ), .ZN(n63) );
  INV_X4 U30 ( .A(n16), .ZN(n64) );
  INV_X4 U32 ( .A(reset), .ZN(n65) );
endmodule


module y_arbiter ( reset, clock, addressY, count2, EOF, MainCount, sig, 
        EOC_Flag, CompStart );
  output [10:0] addressY;
  input [2:0] count2;
  output [4:0] MainCount;
  input reset, clock, EOF, sig, CompStart;
  output EOC_Flag;
  wire   n35, n78, \U3/U3/Z_0 , \U3/U3/Z_1 , \U3/U3/Z_2 , \U3/U3/Z_3 ,
         \U3/U3/Z_4 , \U3/U3/Z_5 , \U3/U3/Z_10 , \U3/U3/DATA3_0 ,
         \U3/U3/DATA3_1 , \U3/U3/DATA3_2 , \U3/U3/DATA3_3 , \U3/U3/DATA3_4 ,
         \U3/U3/DATA3_5 , \U3/U3/DATA3_6 , \U3/U3/DATA3_7 , \U3/U3/DATA3_8 ,
         \U3/U3/DATA3_9 , \U3/U3/DATA3_10 , \U3/U3/DATA2_1 , \U3/U3/DATA2_2 ,
         \U3/U3/DATA2_3 , \U3/U3/DATA2_4 , \U3/U3/DATA2_5 , \U3/U3/DATA2_6 ,
         \U3/U3/DATA2_7 , \U3/U3/DATA2_8 , \U3/U3/DATA2_9 , \U5/Z_0 , \U5/Z_1 ,
         \U5/Z_2 , \U4/DATA2_1 , \U4/DATA2_2 , \U4/DATA2_3 , \U4/DATA2_4 ,
         \add_46/A[0] , \add_46/A[1] , \add_46/A[2] , \sub_98/carry[2] ,
         \sub_98/carry[3] , \sub_98/carry[4] , \sub_98/A[0] , \sub_98/A[1] ,
         \sub_98/A[2] , \sub_98/A[3] , \sub_98/A[4] , \add_79/carry[10] ,
         \add_79/carry[9] , \add_79/carry[8] , \add_79/carry[7] ,
         \add_79/carry[6] , \add_79/carry[5] , \add_79/carry[4] ,
         \add_79/carry[3] , \add_79/carry[2] , \eq_122/B[0] , \eq_122/B[1] ,
         \eq_122/B[2] , n2, n11, n12, n13, n14, n17, n19, n20, n21, n22, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121;
  assign addressY[0] = \U3/U3/DATA3_0 ;
  assign addressY[1] = \U3/U3/DATA3_1 ;
  assign addressY[2] = \U3/U3/DATA3_2 ;
  assign addressY[3] = \U3/U3/DATA3_3 ;
  assign addressY[4] = \U3/U3/DATA3_4 ;
  assign addressY[5] = \U3/U3/DATA3_5 ;
  assign addressY[6] = \U3/U3/DATA3_6 ;
  assign addressY[7] = \U3/U3/DATA3_7 ;
  assign addressY[8] = \U3/U3/DATA3_8 ;
  assign addressY[9] = \U3/U3/DATA3_9 ;
  assign addressY[10] = \U3/U3/DATA3_10 ;
  assign MainCount[0] = \sub_98/A[0] ;
  assign MainCount[1] = \sub_98/A[1] ;
  assign MainCount[2] = \sub_98/A[2] ;
  assign MainCount[3] = \sub_98/A[3] ;
  assign MainCount[4] = \sub_98/A[4] ;
  assign \eq_122/B[0]  = count2[0];
  assign \eq_122/B[1]  = count2[1];
  assign \eq_122/B[2]  = count2[2];

  HA_X1 \add_79/U1_1_1  ( .A(\U3/U3/DATA3_1 ), .B(\U3/U3/DATA3_0 ), .CO(
        \add_79/carry[2] ), .S(\U3/U3/DATA2_1 ) );
  HA_X1 \add_79/U1_1_2  ( .A(\U3/U3/DATA3_2 ), .B(\add_79/carry[2] ), .CO(
        \add_79/carry[3] ), .S(\U3/U3/DATA2_2 ) );
  HA_X1 \add_79/U1_1_3  ( .A(\U3/U3/DATA3_3 ), .B(\add_79/carry[3] ), .CO(
        \add_79/carry[4] ), .S(\U3/U3/DATA2_3 ) );
  HA_X1 \add_79/U1_1_4  ( .A(\U3/U3/DATA3_4 ), .B(\add_79/carry[4] ), .CO(
        \add_79/carry[5] ), .S(\U3/U3/DATA2_4 ) );
  HA_X1 \add_79/U1_1_5  ( .A(\U3/U3/DATA3_5 ), .B(\add_79/carry[5] ), .CO(
        \add_79/carry[6] ), .S(\U3/U3/DATA2_5 ) );
  HA_X1 \add_79/U1_1_6  ( .A(\U3/U3/DATA3_6 ), .B(\add_79/carry[6] ), .CO(
        \add_79/carry[7] ), .S(\U3/U3/DATA2_6 ) );
  HA_X1 \add_79/U1_1_7  ( .A(\U3/U3/DATA3_7 ), .B(\add_79/carry[7] ), .CO(
        \add_79/carry[8] ), .S(\U3/U3/DATA2_7 ) );
  HA_X1 \add_79/U1_1_8  ( .A(\U3/U3/DATA3_8 ), .B(\add_79/carry[8] ), .CO(
        \add_79/carry[9] ), .S(\U3/U3/DATA2_8 ) );
  HA_X1 \add_79/U1_1_9  ( .A(\U3/U3/DATA3_9 ), .B(\add_79/carry[9] ), .CO(
        \add_79/carry[10] ), .S(\U3/U3/DATA2_9 ) );
  XNOR2_X2 \sub_98/U1_A_1  ( .A(\sub_98/A[1] ), .B(\sub_98/A[0] ), .ZN(
        \U4/DATA2_1 ) );
  XNOR2_X2 \sub_98/U1_A_2  ( .A(\sub_98/A[2] ), .B(\sub_98/carry[2] ), .ZN(
        \U4/DATA2_2 ) );
  OR2_X1 \sub_98/U1_B_2  ( .A1(\sub_98/A[2] ), .A2(\sub_98/carry[2] ), .ZN(
        \sub_98/carry[3] ) );
  XNOR2_X2 \sub_98/U1_A_3  ( .A(\sub_98/A[3] ), .B(\sub_98/carry[3] ), .ZN(
        \U4/DATA2_3 ) );
  OR2_X1 \sub_98/U1_B_3  ( .A1(\sub_98/A[3] ), .A2(\sub_98/carry[3] ), .ZN(
        \sub_98/carry[4] ) );
  XNOR2_X2 \sub_98/U1_A_4  ( .A(\sub_98/A[4] ), .B(\sub_98/carry[4] ), .ZN(
        \U4/DATA2_4 ) );
  DFF_X1 \MainCount_reg[0]  ( .D(n67), .CK(clock), .Q(\sub_98/A[0] ), .QN(n22)
         );
  SDFF_X1 NewFlag_reg ( .D(n37), .SI(1'b0), .SE(n121), .CK(clock), .Q(n35) );
  DFF_X1 HoldFlag_reg ( .D(n62), .CK(clock), .Q(n78), .QN(n14) );
  DFF_X1 \count_reg[0]  ( .D(\U5/Z_0 ), .CK(clock), .Q(\add_46/A[0] ) );
  DFF_X1 \count_reg[1]  ( .D(\U5/Z_1 ), .CK(clock), .Q(\add_46/A[1] ), .QN(n11) );
  DFF_X1 \count_reg[2]  ( .D(\U5/Z_2 ), .CK(clock), .Q(\add_46/A[2] ), .QN(n2)
         );
  DFF_X1 \addressY_reg[0]  ( .D(\U3/U3/Z_0 ), .CK(clock), .Q(\U3/U3/DATA3_0 ), 
        .QN(n13) );
  DFF_X1 \addressY_reg[1]  ( .D(\U3/U3/Z_1 ), .CK(clock), .Q(\U3/U3/DATA3_1 )
         );
  DFF_X1 \addressY_reg[2]  ( .D(\U3/U3/Z_2 ), .CK(clock), .Q(\U3/U3/DATA3_2 )
         );
  DFF_X1 \addressY_reg[3]  ( .D(\U3/U3/Z_3 ), .CK(clock), .Q(\U3/U3/DATA3_3 )
         );
  DFF_X1 \addressY_reg[4]  ( .D(\U3/U3/Z_4 ), .CK(clock), .Q(\U3/U3/DATA3_4 )
         );
  DFF_X1 \addressY_reg[5]  ( .D(\U3/U3/Z_5 ), .CK(clock), .Q(\U3/U3/DATA3_5 )
         );
  DFF_X1 \addressY_reg[6]  ( .D(n111), .CK(clock), .Q(\U3/U3/DATA3_6 ) );
  DFF_X1 \addressY_reg[7]  ( .D(n112), .CK(clock), .Q(\U3/U3/DATA3_7 ) );
  DFF_X1 \addressY_reg[8]  ( .D(n113), .CK(clock), .Q(\U3/U3/DATA3_8 ) );
  DFF_X1 \addressY_reg[9]  ( .D(n114), .CK(clock), .Q(\U3/U3/DATA3_9 ) );
  DFF_X1 \MainCount_reg[2]  ( .D(n64), .CK(clock), .Q(\sub_98/A[2] ), .QN(n20)
         );
  DFF_X1 \MainCount_reg[3]  ( .D(n63), .CK(clock), .Q(\sub_98/A[3] ), .QN(n19)
         );
  DFF_X1 \MainCount_reg[4]  ( .D(n66), .CK(clock), .Q(\sub_98/A[4] ), .QN(n17)
         );
  NAND4_X2 U5 ( .A1(n28), .A2(n26), .A3(n119), .A4(n120), .ZN(n27) );
  NAND2_X2 U6 ( .A1(n78), .A2(n29), .ZN(n28) );
  NAND2_X2 U7 ( .A1(n30), .A2(n29), .ZN(n26) );
  NAND2_X2 U9 ( .A1(\U4/DATA2_3 ), .A2(n34), .ZN(n33) );
  NAND2_X2 U11 ( .A1(\U4/DATA2_2 ), .A2(n34), .ZN(n36) );
  NAND2_X2 U13 ( .A1(\U4/DATA2_1 ), .A2(n34), .ZN(n38) );
  NAND2_X2 U15 ( .A1(\U4/DATA2_4 ), .A2(n34), .ZN(n39) );
  OAI22_X2 U16 ( .A1(n32), .A2(n22), .B1(\sub_98/A[0] ), .B2(n108), .ZN(n67)
         );
  NAND2_X2 U17 ( .A1(n37), .A2(n108), .ZN(n32) );
  NOR3_X2 U18 ( .A1(n35), .A2(n121), .A3(n117), .ZN(n34) );
  NAND4_X2 U20 ( .A1(n118), .A2(\add_46/A[1] ), .A3(\add_46/A[0] ), .A4(n2), 
        .ZN(n41) );
  NOR2_X2 U22 ( .A1(n43), .A2(n42), .ZN(\U5/Z_1 ) );
  XNOR2_X2 U23 ( .A(\add_46/A[0] ), .B(\add_46/A[1] ), .ZN(n43) );
  NOR2_X2 U24 ( .A1(n42), .A2(\add_46/A[0] ), .ZN(\U5/Z_0 ) );
  NAND4_X2 U25 ( .A1(n31), .A2(n119), .A3(n14), .A4(n120), .ZN(n42) );
  NAND2_X2 U30 ( .A1(n49), .A2(n30), .ZN(\U3/U3/Z_5 ) );
  NAND2_X2 U32 ( .A1(n50), .A2(n30), .ZN(\U3/U3/Z_4 ) );
  NAND2_X2 U34 ( .A1(n51), .A2(n30), .ZN(\U3/U3/Z_3 ) );
  NAND2_X2 U36 ( .A1(n52), .A2(n30), .ZN(\U3/U3/Z_2 ) );
  NAND3_X2 U39 ( .A1(n116), .A2(n12), .A3(\add_79/carry[10] ), .ZN(n53) );
  NAND2_X2 U41 ( .A1(n56), .A2(n30), .ZN(\U3/U3/Z_1 ) );
  OAI221_X2 U43 ( .B1(n110), .B2(n13), .C1(\U3/U3/DATA3_0 ), .C2(n55), .A(n30), 
        .ZN(\U3/U3/Z_0 ) );
  NAND2_X2 U44 ( .A1(n57), .A2(n30), .ZN(n55) );
  NOR3_X2 U46 ( .A1(EOF), .A2(n78), .A3(n31), .ZN(n57) );
  NAND3_X2 U47 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n31) );
  XNOR2_X2 U48 ( .A(\add_46/A[2] ), .B(\eq_122/B[2] ), .ZN(n60) );
  XNOR2_X2 U49 ( .A(\add_46/A[0] ), .B(\eq_122/B[0] ), .ZN(n59) );
  XNOR2_X2 U50 ( .A(\add_46/A[1] ), .B(\eq_122/B[1] ), .ZN(n58) );
  NOR2_X2 U52 ( .A1(reset), .A2(EOC_Flag), .ZN(n37) );
  AND4_X2 U53 ( .A1(n22), .A2(n21), .A3(sig), .A4(n61), .ZN(EOC_Flag) );
  NOR3_X2 U54 ( .A1(\sub_98/A[2] ), .A2(\sub_98/A[4] ), .A3(\sub_98/A[3] ), 
        .ZN(n61) );
  OR2_X1 U69 ( .A1(n121), .A2(n31), .ZN(n29) );
  DFF_X2 \MainCount_reg[1]  ( .D(n65), .CK(clock), .Q(\sub_98/A[1] ), .QN(n21)
         );
  DFF_X2 \addressY_reg[10]  ( .D(\U3/U3/Z_10 ), .CK(clock), .Q(
        \U3/U3/DATA3_10 ), .QN(n12) );
  NAND2_X2 U4 ( .A1(n21), .A2(n22), .ZN(\sub_98/carry[2] ) );
  INV_X4 U8 ( .A(n55), .ZN(n116) );
  NOR2_X2 U10 ( .A1(n115), .A2(n57), .ZN(n45) );
  AOI211_X1 U12 ( .C1(sig), .C2(n78), .A(CompStart), .B(n117), .ZN(n30) );
  AOI22_X2 U14 ( .A1(\U3/U3/DATA3_5 ), .A2(n45), .B1(\U3/U3/DATA2_5 ), .B2(
        n116), .ZN(n49) );
  AOI22_X2 U19 ( .A1(\U3/U3/DATA3_4 ), .A2(n45), .B1(\U3/U3/DATA2_4 ), .B2(
        n116), .ZN(n50) );
  AOI22_X2 U21 ( .A1(\U3/U3/DATA3_3 ), .A2(n45), .B1(\U3/U3/DATA2_3 ), .B2(
        n116), .ZN(n51) );
  AOI22_X2 U26 ( .A1(\U3/U3/DATA3_2 ), .A2(n45), .B1(\U3/U3/DATA2_2 ), .B2(
        n116), .ZN(n52) );
  AOI22_X2 U27 ( .A1(\U3/U3/DATA3_1 ), .A2(n45), .B1(\U3/U3/DATA2_1 ), .B2(
        n116), .ZN(n56) );
  OAI21_X2 U28 ( .B1(n109), .B2(n12), .A(n53), .ZN(\U3/U3/Z_10 ) );
  OAI21_X2 U29 ( .B1(n55), .B2(\add_79/carry[10] ), .A(n110), .ZN(n54) );
  AOI22_X2 U31 ( .A1(\U3/U3/DATA3_9 ), .A2(n45), .B1(\U3/U3/DATA2_9 ), .B2(
        n116), .ZN(n44) );
  AOI22_X2 U33 ( .A1(\U3/U3/DATA3_8 ), .A2(n45), .B1(\U3/U3/DATA2_8 ), .B2(
        n116), .ZN(n46) );
  AOI22_X2 U35 ( .A1(\U3/U3/DATA3_7 ), .A2(n45), .B1(\U3/U3/DATA2_7 ), .B2(
        n116), .ZN(n47) );
  AOI22_X2 U37 ( .A1(\U3/U3/DATA3_6 ), .A2(n45), .B1(\U3/U3/DATA2_6 ), .B2(
        n116), .ZN(n48) );
  OAI211_X2 U38 ( .C1(n32), .C2(n17), .A(n39), .B(n37), .ZN(n66) );
  OAI211_X2 U40 ( .C1(n32), .C2(n20), .A(n36), .B(n37), .ZN(n64) );
  OAI21_X2 U42 ( .B1(n32), .B2(n21), .A(n38), .ZN(n65) );
  OAI21_X2 U45 ( .B1(n32), .B2(n19), .A(n33), .ZN(n63) );
  OAI21_X2 U51 ( .B1(n14), .B2(n26), .A(n27), .ZN(n62) );
  OAI21_X2 U55 ( .B1(n40), .B2(n2), .A(n41), .ZN(\U5/Z_2 ) );
  AOI21_X2 U56 ( .B1(n118), .B2(n11), .A(\U5/Z_0 ), .ZN(n40) );
  INV_X4 U57 ( .A(n34), .ZN(n108) );
  INV_X4 U58 ( .A(n54), .ZN(n109) );
  INV_X4 U59 ( .A(n45), .ZN(n110) );
  INV_X4 U60 ( .A(n48), .ZN(n111) );
  INV_X4 U61 ( .A(n47), .ZN(n112) );
  INV_X4 U62 ( .A(n46), .ZN(n113) );
  INV_X4 U63 ( .A(n44), .ZN(n114) );
  INV_X4 U64 ( .A(n30), .ZN(n115) );
  INV_X4 U65 ( .A(n37), .ZN(n117) );
  INV_X4 U66 ( .A(n42), .ZN(n118) );
  INV_X4 U67 ( .A(CompStart), .ZN(n119) );
  INV_X4 U68 ( .A(reset), .ZN(n120) );
  INV_X4 U70 ( .A(EOF), .ZN(n121) );
endmodule


module decoder ( clock, reset, data, Diagonal, Element, ElementAddr, EOF, sig, 
        CompStart );
  input [255:0] data;
  output [47:0] Diagonal;
  output [48:0] Element;
  output [10:0] ElementAddr;
  input clock, reset, EOF, sig, CompStart;
  wire   \U3/U5/DATA3_0 , \U3/U5/DATA3_1 , \U3/U5/DATA3_2 , \U3/U5/DATA3_3 ,
         \U3/U5/DATA2_0 , \U3/U5/DATA2_1 , \U3/U5/DATA2_2 , \U3/U5/DATA2_3 ,
         \U3/U5/DATA1_0 , \U3/U5/DATA1_1 , \U3/U5/DATA1_2 , \U3/U5/DATA1_3 ,
         \U27/DATA2_0 , \U27/DATA2_1 , \U27/DATA2_2 , \U27/DATA2_3 ,
         \U27/DATA2_4 , \U27/DATA2_5 , \U27/DATA2_6 , \U27/DATA2_7 ,
         \U27/DATA2_8 , \U27/DATA2_9 , \U27/DATA2_10 , \U27/DATA2_11 ,
         \U27/DATA2_12 , \U27/DATA2_13 , \U27/DATA2_14 , \U27/DATA2_15 ,
         \U27/DATA2_16 , \U27/DATA2_17 , \U27/DATA2_18 , \U27/DATA2_19 ,
         \U27/DATA2_20 , \U27/DATA2_21 , \U27/DATA2_22 , \U27/DATA2_23 ,
         \U27/DATA2_24 , \U27/DATA2_25 , \U27/DATA2_26 , \U27/DATA2_27 ,
         \U27/DATA2_28 , \U27/DATA2_29 , \U27/DATA2_30 , \U27/DATA2_31 ,
         \U27/DATA2_32 , \U27/DATA2_33 , \U27/DATA2_34 , \U27/DATA2_35 ,
         \U27/DATA2_36 , \U27/DATA2_37 , \U27/DATA2_38 , \U27/DATA2_39 ,
         \U27/DATA2_40 , \U27/DATA2_41 , \U27/DATA2_42 , \U27/DATA2_43 ,
         \U27/DATA2_44 , \U27/DATA2_45 , \U27/DATA2_46 , \U27/DATA2_47 ,
         \U27/DATA1_0 , \U27/DATA1_1 , \U27/DATA1_2 , \U27/DATA1_3 ,
         \U27/DATA1_4 , \U27/DATA1_5 , \U27/DATA1_6 , \U27/DATA1_7 ,
         \U27/DATA1_8 , \U27/DATA1_9 , \U27/DATA1_10 , \U27/DATA1_11 ,
         \U27/DATA1_12 , \U27/DATA1_13 , \U27/DATA1_14 , \U27/DATA1_15 ,
         \U27/DATA1_16 , \U27/DATA1_17 , \U27/DATA1_18 , \U27/DATA1_19 ,
         \U27/DATA1_20 , \U27/DATA1_21 , \U27/DATA1_22 , \U27/DATA1_23 ,
         \U27/DATA1_24 , \U27/DATA1_25 , \U27/DATA1_26 , \U27/DATA1_27 ,
         \U27/DATA1_28 , \U27/DATA1_29 , \U27/DATA1_30 , \U27/DATA1_31 ,
         \U27/DATA1_32 , \U27/DATA1_33 , \U27/DATA1_34 , \U27/DATA1_35 ,
         \U27/DATA1_36 , \U27/DATA1_37 , \U27/DATA1_38 , \U27/DATA1_39 ,
         \U27/DATA1_40 , \U27/DATA1_41 , \U27/DATA1_42 , \U27/DATA1_43 ,
         \U27/DATA1_44 , \U27/DATA1_45 , \U27/DATA1_46 , \U27/DATA1_47 ,
         \U26/DATA2_0 , \U26/DATA2_1 , \U26/DATA2_2 , \U26/DATA2_3 ,
         \U26/DATA2_4 , \U26/DATA2_5 , \U26/DATA2_6 , \U26/DATA2_7 ,
         \U26/DATA1_0 , \U26/DATA1_1 , \U26/DATA1_2 , \U26/DATA1_3 ,
         \U26/DATA1_4 , \U26/DATA1_5 , \U26/DATA1_6 , \U26/DATA1_7 ,
         \U24/DATA1_0 , \U24/DATA1_1 , \U24/DATA1_2 , \U24/DATA1_3 ,
         \U24/DATA1_4 , \U24/DATA1_5 , \U24/DATA1_6 , \U24/DATA1_7 ,
         \U24/DATA1_8 , \U24/DATA1_9 , \U24/DATA1_10 , \U24/DATA1_11 ,
         \U24/DATA1_12 , \U24/DATA1_13 , \U24/DATA1_14 , \U24/DATA1_15 ,
         \U24/DATA1_16 , \U24/DATA1_17 , \U24/DATA1_18 , \U24/DATA1_19 ,
         \U24/DATA1_20 , \U24/DATA1_21 , \U24/DATA1_22 , \U24/DATA1_23 ,
         \U24/DATA1_24 , \U24/DATA1_25 , \U24/DATA1_26 , \U24/DATA1_27 ,
         \U24/DATA1_28 , \U24/DATA1_29 , \U24/DATA1_30 , \U24/DATA1_31 ,
         \U24/DATA1_32 , \U24/DATA1_33 , \U24/DATA1_34 , \U24/DATA1_35 ,
         \U24/DATA1_36 , \U24/DATA1_37 , \U24/DATA1_38 , \U24/DATA1_39 ,
         \U24/DATA1_40 , \U24/DATA1_41 , \U24/DATA1_42 , \U24/DATA1_43 ,
         \U24/DATA1_44 , \U24/DATA1_45 , \U24/DATA1_46 , \U24/DATA1_47 ,
         \U23/DATA1_0 , \U23/DATA1_1 , \U23/DATA1_2 , \U23/DATA1_3 ,
         \U23/DATA1_4 , \U23/DATA1_5 , \U23/DATA1_6 , \U23/DATA1_7 ,
         \U21/DATA1_0 , \U21/DATA1_1 , \U21/DATA1_2 , \U21/DATA1_3 ,
         \U21/DATA1_4 , \U21/DATA1_5 , \U21/DATA1_6 , \U21/DATA1_7 ,
         \U21/DATA1_8 , \U21/DATA1_9 , \U21/DATA1_10 , \U21/DATA1_11 ,
         \U21/DATA1_12 , \U21/DATA1_13 , \U21/DATA1_14 , \U21/DATA1_15 ,
         \U21/DATA1_16 , \U21/DATA1_17 , \U21/DATA1_18 , \U21/DATA1_19 ,
         \U21/DATA1_20 , \U21/DATA1_21 , \U21/DATA1_22 , \U21/DATA1_23 ,
         \U21/DATA1_24 , \U21/DATA1_25 , \U21/DATA1_26 , \U21/DATA1_27 ,
         \U21/DATA1_28 , \U21/DATA1_29 , \U21/DATA1_30 , \U21/DATA1_31 ,
         \U21/DATA1_32 , \U21/DATA1_33 , \U21/DATA1_34 , \U21/DATA1_35 ,
         \U21/DATA1_36 , \U21/DATA1_37 , \U21/DATA1_38 , \U21/DATA1_39 ,
         \U21/DATA1_40 , \U21/DATA1_41 , \U21/DATA1_42 , \U21/DATA1_43 ,
         \U21/DATA1_44 , \U21/DATA1_45 , \U21/DATA1_46 , \U21/DATA1_47 ,
         \U20/DATA1_0 , \U20/DATA1_1 , \U20/DATA1_2 , \U20/DATA1_3 ,
         \U20/DATA1_4 , \U20/DATA1_5 , \U20/DATA1_6 , \U20/DATA1_7 ,
         \U20/DATA1_8 , \U20/DATA1_9 , \U20/DATA1_10 , \U4/DATA4_3 ,
         \r412/A[0] , \r412/A[1] , \r389/A[0] , \r389/A[1] , \r389/A[2] ,
         \r389/A[3] , n16, n120, n121, n122, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996;
  assign \U3/U5/DATA3_0  = data[248];
  assign \U3/U5/DATA3_1  = data[249];
  assign \U3/U5/DATA3_2  = data[250];
  assign \U3/U5/DATA3_3  = data[251];
  assign \U3/U5/DATA2_0  = data[184];
  assign \U3/U5/DATA2_1  = data[185];
  assign \U3/U5/DATA2_2  = data[186];
  assign \U3/U5/DATA2_3  = data[187];
  assign \U3/U5/DATA1_0  = data[120];
  assign \U3/U5/DATA1_1  = data[121];
  assign \U3/U5/DATA1_2  = data[122];
  assign \U3/U5/DATA1_3  = data[123];
  assign \U27/DATA2_0  = data[192];
  assign \U27/DATA2_1  = data[193];
  assign \U27/DATA2_2  = data[194];
  assign \U27/DATA2_3  = data[195];
  assign \U27/DATA2_4  = data[196];
  assign \U27/DATA2_5  = data[197];
  assign \U27/DATA2_6  = data[198];
  assign \U27/DATA2_7  = data[199];
  assign \U27/DATA2_8  = data[200];
  assign \U27/DATA2_9  = data[201];
  assign \U27/DATA2_10  = data[202];
  assign \U27/DATA2_11  = data[203];
  assign \U27/DATA2_12  = data[204];
  assign \U27/DATA2_13  = data[205];
  assign \U27/DATA2_14  = data[206];
  assign \U27/DATA2_15  = data[207];
  assign \U27/DATA2_16  = data[208];
  assign \U27/DATA2_17  = data[209];
  assign \U27/DATA2_18  = data[210];
  assign \U27/DATA2_19  = data[211];
  assign \U27/DATA2_20  = data[212];
  assign \U27/DATA2_21  = data[213];
  assign \U27/DATA2_22  = data[214];
  assign \U27/DATA2_23  = data[215];
  assign \U27/DATA2_24  = data[216];
  assign \U27/DATA2_25  = data[217];
  assign \U27/DATA2_26  = data[218];
  assign \U27/DATA2_27  = data[219];
  assign \U27/DATA2_28  = data[220];
  assign \U27/DATA2_29  = data[221];
  assign \U27/DATA2_30  = data[222];
  assign \U27/DATA2_31  = data[223];
  assign \U27/DATA2_32  = data[224];
  assign \U27/DATA2_33  = data[225];
  assign \U27/DATA2_34  = data[226];
  assign \U27/DATA2_35  = data[227];
  assign \U27/DATA2_36  = data[228];
  assign \U27/DATA2_37  = data[229];
  assign \U27/DATA2_38  = data[230];
  assign \U27/DATA2_39  = data[231];
  assign \U27/DATA2_40  = data[232];
  assign \U27/DATA2_41  = data[233];
  assign \U27/DATA2_42  = data[234];
  assign \U27/DATA2_43  = data[235];
  assign \U27/DATA2_44  = data[236];
  assign \U27/DATA2_45  = data[237];
  assign \U27/DATA2_46  = data[238];
  assign \U27/DATA2_47  = data[239];
  assign \U27/DATA1_0  = data[128];
  assign \U27/DATA1_1  = data[129];
  assign \U27/DATA1_2  = data[130];
  assign \U27/DATA1_3  = data[131];
  assign \U27/DATA1_4  = data[132];
  assign \U27/DATA1_5  = data[133];
  assign \U27/DATA1_6  = data[134];
  assign \U27/DATA1_7  = data[135];
  assign \U27/DATA1_8  = data[136];
  assign \U27/DATA1_9  = data[137];
  assign \U27/DATA1_10  = data[138];
  assign \U27/DATA1_11  = data[139];
  assign \U27/DATA1_12  = data[140];
  assign \U27/DATA1_13  = data[141];
  assign \U27/DATA1_14  = data[142];
  assign \U27/DATA1_15  = data[143];
  assign \U27/DATA1_16  = data[144];
  assign \U27/DATA1_17  = data[145];
  assign \U27/DATA1_18  = data[146];
  assign \U27/DATA1_19  = data[147];
  assign \U27/DATA1_20  = data[148];
  assign \U27/DATA1_21  = data[149];
  assign \U27/DATA1_22  = data[150];
  assign \U27/DATA1_23  = data[151];
  assign \U27/DATA1_24  = data[152];
  assign \U27/DATA1_25  = data[153];
  assign \U27/DATA1_26  = data[154];
  assign \U27/DATA1_27  = data[155];
  assign \U27/DATA1_28  = data[156];
  assign \U27/DATA1_29  = data[157];
  assign \U27/DATA1_30  = data[158];
  assign \U27/DATA1_31  = data[159];
  assign \U27/DATA1_32  = data[160];
  assign \U27/DATA1_33  = data[161];
  assign \U27/DATA1_34  = data[162];
  assign \U27/DATA1_35  = data[163];
  assign \U27/DATA1_36  = data[164];
  assign \U27/DATA1_37  = data[165];
  assign \U27/DATA1_38  = data[166];
  assign \U27/DATA1_39  = data[167];
  assign \U27/DATA1_40  = data[168];
  assign \U27/DATA1_41  = data[169];
  assign \U27/DATA1_42  = data[170];
  assign \U27/DATA1_43  = data[171];
  assign \U27/DATA1_44  = data[172];
  assign \U27/DATA1_45  = data[173];
  assign \U27/DATA1_46  = data[174];
  assign \U27/DATA1_47  = data[175];
  assign \U26/DATA2_0  = data[240];
  assign \U26/DATA2_1  = data[241];
  assign \U26/DATA2_2  = data[242];
  assign \U26/DATA2_3  = data[243];
  assign \U26/DATA2_4  = data[244];
  assign \U26/DATA2_5  = data[245];
  assign \U26/DATA2_6  = data[246];
  assign \U26/DATA2_7  = data[247];
  assign \U26/DATA1_0  = data[176];
  assign \U26/DATA1_1  = data[177];
  assign \U26/DATA1_2  = data[178];
  assign \U26/DATA1_3  = data[179];
  assign \U26/DATA1_4  = data[180];
  assign \U26/DATA1_5  = data[181];
  assign \U26/DATA1_6  = data[182];
  assign \U26/DATA1_7  = data[183];
  assign \U24/DATA1_0  = data[64];
  assign \U24/DATA1_1  = data[65];
  assign \U24/DATA1_2  = data[66];
  assign \U24/DATA1_3  = data[67];
  assign \U24/DATA1_4  = data[68];
  assign \U24/DATA1_5  = data[69];
  assign \U24/DATA1_6  = data[70];
  assign \U24/DATA1_7  = data[71];
  assign \U24/DATA1_8  = data[72];
  assign \U24/DATA1_9  = data[73];
  assign \U24/DATA1_10  = data[74];
  assign \U24/DATA1_11  = data[75];
  assign \U24/DATA1_12  = data[76];
  assign \U24/DATA1_13  = data[77];
  assign \U24/DATA1_14  = data[78];
  assign \U24/DATA1_15  = data[79];
  assign \U24/DATA1_16  = data[80];
  assign \U24/DATA1_17  = data[81];
  assign \U24/DATA1_18  = data[82];
  assign \U24/DATA1_19  = data[83];
  assign \U24/DATA1_20  = data[84];
  assign \U24/DATA1_21  = data[85];
  assign \U24/DATA1_22  = data[86];
  assign \U24/DATA1_23  = data[87];
  assign \U24/DATA1_24  = data[88];
  assign \U24/DATA1_25  = data[89];
  assign \U24/DATA1_26  = data[90];
  assign \U24/DATA1_27  = data[91];
  assign \U24/DATA1_28  = data[92];
  assign \U24/DATA1_29  = data[93];
  assign \U24/DATA1_30  = data[94];
  assign \U24/DATA1_31  = data[95];
  assign \U24/DATA1_32  = data[96];
  assign \U24/DATA1_33  = data[97];
  assign \U24/DATA1_34  = data[98];
  assign \U24/DATA1_35  = data[99];
  assign \U24/DATA1_36  = data[100];
  assign \U24/DATA1_37  = data[101];
  assign \U24/DATA1_38  = data[102];
  assign \U24/DATA1_39  = data[103];
  assign \U24/DATA1_40  = data[104];
  assign \U24/DATA1_41  = data[105];
  assign \U24/DATA1_42  = data[106];
  assign \U24/DATA1_43  = data[107];
  assign \U24/DATA1_44  = data[108];
  assign \U24/DATA1_45  = data[109];
  assign \U24/DATA1_46  = data[110];
  assign \U24/DATA1_47  = data[111];
  assign \U23/DATA1_0  = data[112];
  assign \U23/DATA1_1  = data[113];
  assign \U23/DATA1_2  = data[114];
  assign \U23/DATA1_3  = data[115];
  assign \U23/DATA1_4  = data[116];
  assign \U23/DATA1_5  = data[117];
  assign \U23/DATA1_6  = data[118];
  assign \U23/DATA1_7  = data[119];
  assign \U21/DATA1_0  = data[0];
  assign \U21/DATA1_1  = data[1];
  assign \U21/DATA1_2  = data[2];
  assign \U21/DATA1_3  = data[3];
  assign \U21/DATA1_4  = data[4];
  assign \U21/DATA1_5  = data[5];
  assign \U21/DATA1_6  = data[6];
  assign \U21/DATA1_7  = data[7];
  assign \U21/DATA1_8  = data[8];
  assign \U21/DATA1_9  = data[9];
  assign \U21/DATA1_10  = data[10];
  assign \U21/DATA1_11  = data[11];
  assign \U21/DATA1_12  = data[12];
  assign \U21/DATA1_13  = data[13];
  assign \U21/DATA1_14  = data[14];
  assign \U21/DATA1_15  = data[15];
  assign \U21/DATA1_16  = data[16];
  assign \U21/DATA1_17  = data[17];
  assign \U21/DATA1_18  = data[18];
  assign \U21/DATA1_19  = data[19];
  assign \U21/DATA1_20  = data[20];
  assign \U21/DATA1_21  = data[21];
  assign \U21/DATA1_22  = data[22];
  assign \U21/DATA1_23  = data[23];
  assign \U21/DATA1_24  = data[24];
  assign \U21/DATA1_25  = data[25];
  assign \U21/DATA1_26  = data[26];
  assign \U21/DATA1_27  = data[27];
  assign \U21/DATA1_28  = data[28];
  assign \U21/DATA1_29  = data[29];
  assign \U21/DATA1_30  = data[30];
  assign \U21/DATA1_31  = data[31];
  assign \U21/DATA1_32  = data[32];
  assign \U21/DATA1_33  = data[33];
  assign \U21/DATA1_34  = data[34];
  assign \U21/DATA1_35  = data[35];
  assign \U21/DATA1_36  = data[36];
  assign \U21/DATA1_37  = data[37];
  assign \U21/DATA1_38  = data[38];
  assign \U21/DATA1_39  = data[39];
  assign \U21/DATA1_40  = data[40];
  assign \U21/DATA1_41  = data[41];
  assign \U21/DATA1_42  = data[42];
  assign \U21/DATA1_43  = data[43];
  assign \U21/DATA1_44  = data[44];
  assign \U21/DATA1_45  = data[45];
  assign \U21/DATA1_46  = data[46];
  assign \U21/DATA1_47  = data[47];
  assign \U20/DATA1_0  = data[48];
  assign \U20/DATA1_1  = data[49];
  assign \U20/DATA1_2  = data[50];
  assign \U20/DATA1_3  = data[51];
  assign \U20/DATA1_4  = data[52];
  assign \U20/DATA1_5  = data[53];
  assign \U20/DATA1_6  = data[54];
  assign \U20/DATA1_7  = data[55];
  assign \U20/DATA1_8  = data[56];
  assign \U20/DATA1_9  = data[57];
  assign \U20/DATA1_10  = data[58];
  assign \U4/DATA4_3  = data[59];

  DFF_X1 \Pos_reg[0]  ( .D(n477), .CK(clock), .Q(\r412/A[0] ), .QN(n16) );
  DFF_X1 \NZE_reg[3]  ( .D(n481), .CK(clock), .Q(\r389/A[3] ) );
  DFF_X1 \Pos_reg[1]  ( .D(n476), .CK(clock), .Q(\r412/A[1] ) );
  DFF_X1 \Diagonal_reg[47]  ( .D(n369), .CK(clock), .Q(Diagonal[47]) );
  DFF_X1 \Diagonal_reg[46]  ( .D(n370), .CK(clock), .Q(Diagonal[46]) );
  DFF_X1 \Diagonal_reg[45]  ( .D(n371), .CK(clock), .Q(Diagonal[45]) );
  DFF_X1 \Diagonal_reg[44]  ( .D(n372), .CK(clock), .Q(Diagonal[44]) );
  DFF_X1 \Diagonal_reg[43]  ( .D(n373), .CK(clock), .Q(Diagonal[43]) );
  DFF_X1 \Diagonal_reg[42]  ( .D(n374), .CK(clock), .Q(Diagonal[42]) );
  DFF_X1 \Diagonal_reg[41]  ( .D(n375), .CK(clock), .Q(Diagonal[41]) );
  DFF_X1 \Diagonal_reg[40]  ( .D(n376), .CK(clock), .Q(Diagonal[40]) );
  DFF_X1 \Diagonal_reg[39]  ( .D(n377), .CK(clock), .Q(Diagonal[39]) );
  DFF_X1 \Diagonal_reg[38]  ( .D(n378), .CK(clock), .Q(Diagonal[38]) );
  DFF_X1 \Diagonal_reg[37]  ( .D(n379), .CK(clock), .Q(Diagonal[37]) );
  DFF_X1 \Diagonal_reg[36]  ( .D(n380), .CK(clock), .Q(Diagonal[36]) );
  DFF_X1 \Diagonal_reg[35]  ( .D(n381), .CK(clock), .Q(Diagonal[35]) );
  DFF_X1 \Diagonal_reg[34]  ( .D(n382), .CK(clock), .Q(Diagonal[34]) );
  DFF_X1 \Diagonal_reg[33]  ( .D(n383), .CK(clock), .Q(Diagonal[33]) );
  DFF_X1 \Diagonal_reg[32]  ( .D(n384), .CK(clock), .Q(Diagonal[32]) );
  DFF_X1 \Diagonal_reg[31]  ( .D(n385), .CK(clock), .Q(Diagonal[31]) );
  DFF_X1 \Diagonal_reg[30]  ( .D(n386), .CK(clock), .Q(Diagonal[30]) );
  DFF_X1 \Diagonal_reg[29]  ( .D(n387), .CK(clock), .Q(Diagonal[29]) );
  DFF_X1 \Diagonal_reg[28]  ( .D(n388), .CK(clock), .Q(Diagonal[28]) );
  DFF_X1 \Diagonal_reg[27]  ( .D(n389), .CK(clock), .Q(Diagonal[27]) );
  DFF_X1 \Diagonal_reg[26]  ( .D(n390), .CK(clock), .Q(Diagonal[26]) );
  DFF_X1 \Diagonal_reg[25]  ( .D(n391), .CK(clock), .Q(Diagonal[25]) );
  DFF_X1 \Diagonal_reg[24]  ( .D(n392), .CK(clock), .Q(Diagonal[24]) );
  DFF_X1 \Diagonal_reg[23]  ( .D(n393), .CK(clock), .Q(Diagonal[23]) );
  DFF_X1 \Diagonal_reg[22]  ( .D(n394), .CK(clock), .Q(Diagonal[22]) );
  DFF_X1 \Diagonal_reg[21]  ( .D(n395), .CK(clock), .Q(Diagonal[21]) );
  DFF_X1 \Diagonal_reg[20]  ( .D(n396), .CK(clock), .Q(Diagonal[20]) );
  DFF_X1 \Diagonal_reg[19]  ( .D(n397), .CK(clock), .Q(Diagonal[19]) );
  DFF_X1 \Diagonal_reg[18]  ( .D(n398), .CK(clock), .Q(Diagonal[18]) );
  DFF_X1 \Diagonal_reg[17]  ( .D(n399), .CK(clock), .Q(Diagonal[17]) );
  DFF_X1 \Diagonal_reg[16]  ( .D(n400), .CK(clock), .Q(Diagonal[16]) );
  DFF_X1 \Diagonal_reg[15]  ( .D(n401), .CK(clock), .Q(Diagonal[15]) );
  DFF_X1 \Diagonal_reg[14]  ( .D(n402), .CK(clock), .Q(Diagonal[14]) );
  DFF_X1 \Diagonal_reg[13]  ( .D(n403), .CK(clock), .Q(Diagonal[13]) );
  DFF_X1 \Diagonal_reg[12]  ( .D(n404), .CK(clock), .Q(Diagonal[12]) );
  DFF_X1 \Diagonal_reg[11]  ( .D(n405), .CK(clock), .Q(Diagonal[11]) );
  DFF_X1 \Diagonal_reg[10]  ( .D(n406), .CK(clock), .Q(Diagonal[10]) );
  DFF_X1 \Diagonal_reg[9]  ( .D(n407), .CK(clock), .Q(Diagonal[9]) );
  DFF_X1 \Diagonal_reg[8]  ( .D(n408), .CK(clock), .Q(Diagonal[8]) );
  DFF_X1 \Diagonal_reg[7]  ( .D(n409), .CK(clock), .Q(Diagonal[7]) );
  DFF_X1 \Diagonal_reg[6]  ( .D(n410), .CK(clock), .Q(Diagonal[6]) );
  DFF_X1 \Diagonal_reg[5]  ( .D(n411), .CK(clock), .Q(Diagonal[5]) );
  DFF_X1 \Diagonal_reg[4]  ( .D(n412), .CK(clock), .Q(Diagonal[4]) );
  DFF_X1 \Diagonal_reg[3]  ( .D(n413), .CK(clock), .Q(Diagonal[3]) );
  DFF_X1 \Diagonal_reg[2]  ( .D(n414), .CK(clock), .Q(Diagonal[2]) );
  DFF_X1 \Diagonal_reg[1]  ( .D(n415), .CK(clock), .Q(Diagonal[1]) );
  DFF_X1 \Diagonal_reg[0]  ( .D(n416), .CK(clock), .Q(Diagonal[0]) );
  DFF_X1 \NZE_reg[0]  ( .D(n478), .CK(clock), .Q(\r389/A[0] ) );
  DFF_X1 \NZE_reg[1]  ( .D(n479), .CK(clock), .Q(\r389/A[1] ) );
  DFF_X1 \NZE_reg[2]  ( .D(n480), .CK(clock), .Q(\r389/A[2] ) );
  DFF_X1 \ElementAddr_reg[10]  ( .D(n417), .CK(clock), .Q(ElementAddr[10]) );
  DFF_X1 \ElementAddr_reg[9]  ( .D(n418), .CK(clock), .Q(ElementAddr[9]) );
  DFF_X1 \ElementAddr_reg[8]  ( .D(n419), .CK(clock), .Q(ElementAddr[8]) );
  DFF_X1 \ElementAddr_reg[7]  ( .D(n420), .CK(clock), .Q(ElementAddr[7]) );
  DFF_X1 \ElementAddr_reg[6]  ( .D(n421), .CK(clock), .Q(ElementAddr[6]) );
  DFF_X1 \ElementAddr_reg[5]  ( .D(n422), .CK(clock), .Q(ElementAddr[5]) );
  DFF_X1 \ElementAddr_reg[4]  ( .D(n423), .CK(clock), .Q(ElementAddr[4]) );
  DFF_X1 \ElementAddr_reg[3]  ( .D(n424), .CK(clock), .Q(ElementAddr[3]) );
  DFF_X1 \ElementAddr_reg[2]  ( .D(n425), .CK(clock), .Q(ElementAddr[2]) );
  DFF_X1 \ElementAddr_reg[1]  ( .D(n426), .CK(clock), .Q(ElementAddr[1]) );
  DFF_X1 \ElementAddr_reg[0]  ( .D(n427), .CK(clock), .Q(ElementAddr[0]) );
  DFF_X1 \Element_reg[0]  ( .D(n428), .CK(clock), .Q(Element[0]) );
  DFF_X1 \Element_reg[1]  ( .D(n429), .CK(clock), .Q(Element[1]) );
  DFF_X1 \Element_reg[2]  ( .D(n430), .CK(clock), .Q(Element[2]) );
  DFF_X1 \Element_reg[3]  ( .D(n431), .CK(clock), .Q(Element[3]) );
  DFF_X1 \Element_reg[4]  ( .D(n432), .CK(clock), .Q(Element[4]) );
  DFF_X1 \Element_reg[5]  ( .D(n433), .CK(clock), .Q(Element[5]) );
  DFF_X1 \Element_reg[6]  ( .D(n434), .CK(clock), .Q(Element[6]) );
  DFF_X1 \Element_reg[7]  ( .D(n435), .CK(clock), .Q(Element[7]) );
  DFF_X1 \Element_reg[8]  ( .D(n436), .CK(clock), .Q(Element[8]) );
  DFF_X1 \Element_reg[9]  ( .D(n437), .CK(clock), .Q(Element[9]) );
  DFF_X1 \Element_reg[10]  ( .D(n438), .CK(clock), .Q(Element[10]) );
  DFF_X1 \Element_reg[11]  ( .D(n439), .CK(clock), .Q(Element[11]) );
  DFF_X1 \Element_reg[12]  ( .D(n440), .CK(clock), .Q(Element[12]) );
  DFF_X1 \Element_reg[13]  ( .D(n441), .CK(clock), .Q(Element[13]) );
  DFF_X1 \Element_reg[14]  ( .D(n442), .CK(clock), .Q(Element[14]) );
  DFF_X1 \Element_reg[15]  ( .D(n443), .CK(clock), .Q(Element[15]) );
  DFF_X1 \Element_reg[16]  ( .D(n444), .CK(clock), .Q(Element[16]) );
  DFF_X1 \Element_reg[17]  ( .D(n445), .CK(clock), .Q(Element[17]) );
  DFF_X1 \Element_reg[18]  ( .D(n446), .CK(clock), .Q(Element[18]) );
  DFF_X1 \Element_reg[19]  ( .D(n447), .CK(clock), .Q(Element[19]) );
  DFF_X1 \Element_reg[20]  ( .D(n448), .CK(clock), .Q(Element[20]) );
  DFF_X1 \Element_reg[21]  ( .D(n449), .CK(clock), .Q(Element[21]) );
  DFF_X1 \Element_reg[22]  ( .D(n450), .CK(clock), .Q(Element[22]) );
  DFF_X1 \Element_reg[23]  ( .D(n451), .CK(clock), .Q(Element[23]) );
  DFF_X1 \Element_reg[24]  ( .D(n452), .CK(clock), .Q(Element[24]) );
  DFF_X1 \Element_reg[25]  ( .D(n453), .CK(clock), .Q(Element[25]) );
  DFF_X1 \Element_reg[26]  ( .D(n454), .CK(clock), .Q(Element[26]) );
  DFF_X1 \Element_reg[27]  ( .D(n455), .CK(clock), .Q(Element[27]) );
  DFF_X1 \Element_reg[28]  ( .D(n456), .CK(clock), .Q(Element[28]) );
  DFF_X1 \Element_reg[29]  ( .D(n457), .CK(clock), .Q(Element[29]) );
  DFF_X1 \Element_reg[30]  ( .D(n458), .CK(clock), .Q(Element[30]) );
  DFF_X1 \Element_reg[31]  ( .D(n459), .CK(clock), .Q(Element[31]) );
  DFF_X1 \Element_reg[32]  ( .D(n460), .CK(clock), .Q(Element[32]) );
  DFF_X1 \Element_reg[33]  ( .D(n461), .CK(clock), .Q(Element[33]) );
  DFF_X1 \Element_reg[34]  ( .D(n462), .CK(clock), .Q(Element[34]) );
  DFF_X1 \Element_reg[35]  ( .D(n463), .CK(clock), .Q(Element[35]) );
  DFF_X1 \Element_reg[36]  ( .D(n464), .CK(clock), .Q(Element[36]) );
  DFF_X1 \Element_reg[37]  ( .D(n465), .CK(clock), .Q(Element[37]) );
  DFF_X1 \Element_reg[38]  ( .D(n466), .CK(clock), .Q(Element[38]) );
  DFF_X1 \Element_reg[39]  ( .D(n467), .CK(clock), .Q(Element[39]) );
  DFF_X1 \Element_reg[40]  ( .D(n468), .CK(clock), .Q(Element[40]) );
  DFF_X1 \Element_reg[41]  ( .D(n469), .CK(clock), .Q(Element[41]) );
  DFF_X1 \Element_reg[42]  ( .D(n470), .CK(clock), .Q(Element[42]) );
  DFF_X1 \Element_reg[43]  ( .D(n471), .CK(clock), .Q(Element[43]) );
  DFF_X1 \Element_reg[44]  ( .D(n472), .CK(clock), .Q(Element[44]) );
  DFF_X1 \Element_reg[45]  ( .D(n473), .CK(clock), .Q(Element[45]) );
  DFF_X1 \Element_reg[46]  ( .D(n474), .CK(clock), .Q(Element[46]) );
  DFF_X1 \Element_reg[47]  ( .D(n475), .CK(clock), .Q(Element[47]) );
  DFF_X1 \Element_reg[48]  ( .D(n889), .CK(clock), .Q(Element[48]) );
  NAND2_X2 U156 ( .A1(n230), .A2(n231), .ZN(n420) );
  NAND2_X2 U159 ( .A1(n233), .A2(n234), .ZN(n421) );
  NAND2_X2 U162 ( .A1(n235), .A2(n236), .ZN(n422) );
  NAND2_X2 U165 ( .A1(n237), .A2(n238), .ZN(n423) );
  NAND2_X2 U168 ( .A1(n239), .A2(n240), .ZN(n424) );
  NAND2_X2 U171 ( .A1(n241), .A2(n242), .ZN(n425) );
  NAND2_X2 U174 ( .A1(n243), .A2(n244), .ZN(n426) );
  NAND2_X2 U177 ( .A1(n245), .A2(n246), .ZN(n427) );
  NAND2_X2 U324 ( .A1(n346), .A2(n347), .ZN(n219) );
  NOR2_X2 U328 ( .A1(n345), .A2(n885), .ZN(n224) );
  NAND2_X2 U330 ( .A1(n351), .A2(n349), .ZN(n345) );
  OAI22_X2 U333 ( .A1(\r412/A[1] ), .A2(n888), .B1(n353), .B2(n891), .ZN(n476)
         );
  NAND2_X2 U335 ( .A1(n348), .A2(n347), .ZN(n120) );
  XOR2_X2 U342 ( .A(n356), .B(n361), .Z(n358) );
  OAI221_X2 U343 ( .B1(n247), .B2(n362), .C1(n868), .C2(n993), .A(n363), .ZN(
        n481) );
  NAND3_X2 U344 ( .A1(n351), .A2(n892), .A3(\r389/A[3] ), .ZN(n363) );
  NOR2_X2 U345 ( .A1(n364), .A2(reset), .ZN(n351) );
  NAND2_X2 U347 ( .A1(\r412/A[0] ), .A2(\r412/A[1] ), .ZN(n349) );
  XOR2_X2 U348 ( .A(n365), .B(n366), .Z(n362) );
  NOR2_X2 U350 ( .A1(n884), .A2(n883), .ZN(n356) );
  NOR2_X2 U355 ( .A1(n890), .A2(reset), .ZN(n347) );
  NOR2_X2 U356 ( .A1(n892), .A2(\r389/A[3] ), .ZN(n364) );
  NOR2_X2 U357 ( .A1(n893), .A2(\r389/A[2] ), .ZN(n360) );
  NOR2_X2 U358 ( .A1(\r389/A[1] ), .A2(\r389/A[0] ), .ZN(n357) );
  NOR2_X2 U359 ( .A1(n886), .A2(n348), .ZN(n353) );
  NOR2_X2 U360 ( .A1(n16), .A2(\r412/A[1] ), .ZN(n348) );
  NAND2_X2 U361 ( .A1(\r412/A[1] ), .A2(n16), .ZN(n350) );
  NOR2_X2 U362 ( .A1(\r412/A[0] ), .A2(\r412/A[1] ), .ZN(n346) );
  AND2_X1 U482 ( .A1(n356), .A2(n361), .ZN(n366) );
  NOR2_X4 U3 ( .A1(n351), .A2(n347), .ZN(n866) );
  OR2_X4 U4 ( .A1(n350), .A2(n888), .ZN(n867) );
  OR2_X4 U5 ( .A1(n349), .A2(n888), .ZN(n868) );
  INV_X4 U6 ( .A(n232), .ZN(n869) );
  INV_X4 U7 ( .A(n232), .ZN(n870) );
  INV_X4 U8 ( .A(n873), .ZN(n872) );
  INV_X4 U9 ( .A(n875), .ZN(n874) );
  INV_X4 U10 ( .A(n224), .ZN(n875) );
  INV_X4 U11 ( .A(n878), .ZN(n876) );
  INV_X4 U12 ( .A(n878), .ZN(n877) );
  INV_X4 U13 ( .A(n868), .ZN(n880) );
  INV_X4 U14 ( .A(n881), .ZN(n882) );
  INV_X4 U15 ( .A(n219), .ZN(n871) );
  INV_X4 U16 ( .A(n225), .ZN(n873) );
  INV_X4 U17 ( .A(n222), .ZN(n878) );
  INV_X4 U18 ( .A(n867), .ZN(n879) );
  OAI21_X2 U19 ( .B1(n349), .B2(n891), .A(n867), .ZN(n225) );
  AOI222_X1 U20 ( .A1(n886), .A2(\U3/U5/DATA1_2 ), .B1(n348), .B2(
        \U3/U5/DATA2_2 ), .C1(n346), .C2(\U3/U5/DATA3_2 ), .ZN(n361) );
  AOI222_X1 U21 ( .A1(n886), .A2(\U3/U5/DATA1_0 ), .B1(n348), .B2(
        \U3/U5/DATA2_0 ), .C1(n346), .C2(\U3/U5/DATA3_0 ), .ZN(n367) );
  AOI222_X1 U22 ( .A1(n886), .A2(\U3/U5/DATA1_1 ), .B1(n348), .B2(
        \U3/U5/DATA2_1 ), .C1(n346), .C2(\U3/U5/DATA3_1 ), .ZN(n368) );
  AOI222_X1 U23 ( .A1(\U3/U5/DATA3_3 ), .A2(n346), .B1(\U3/U5/DATA2_3 ), .B2(
        n348), .C1(\U3/U5/DATA1_3 ), .C2(n886), .ZN(n365) );
  OAI21_X2 U24 ( .B1(n346), .B2(n885), .A(n347), .ZN(n247) );
  INV_X4 U25 ( .A(n120), .ZN(n881) );
  OAI21_X2 U26 ( .B1(n887), .B2(n345), .A(n219), .ZN(n222) );
  OAI21_X2 U27 ( .B1(n350), .B2(n345), .A(n882), .ZN(n232) );
  AOI22_X2 U28 ( .A1(\U26/DATA1_0 ), .A2(n222), .B1(ElementAddr[0]), .B2(n223), 
        .ZN(n245) );
  AOI222_X1 U29 ( .A1(\U23/DATA1_0 ), .A2(n232), .B1(\U26/DATA2_0 ), .B2(n874), 
        .C1(\U20/DATA1_0 ), .C2(n225), .ZN(n246) );
  AOI22_X2 U30 ( .A1(\U26/DATA1_1 ), .A2(n876), .B1(ElementAddr[1]), .B2(n223), 
        .ZN(n243) );
  AOI222_X1 U31 ( .A1(\U23/DATA1_1 ), .A2(n232), .B1(\U26/DATA2_1 ), .B2(n874), 
        .C1(\U20/DATA1_1 ), .C2(n225), .ZN(n244) );
  AOI22_X2 U32 ( .A1(\U26/DATA1_2 ), .A2(n877), .B1(ElementAddr[2]), .B2(n223), 
        .ZN(n241) );
  AOI222_X1 U33 ( .A1(\U23/DATA1_2 ), .A2(n232), .B1(\U26/DATA2_2 ), .B2(n874), 
        .C1(\U20/DATA1_2 ), .C2(n225), .ZN(n242) );
  AOI22_X2 U34 ( .A1(\U26/DATA1_3 ), .A2(n222), .B1(ElementAddr[3]), .B2(n223), 
        .ZN(n239) );
  AOI222_X1 U35 ( .A1(\U23/DATA1_3 ), .A2(n232), .B1(\U26/DATA2_3 ), .B2(n874), 
        .C1(\U20/DATA1_3 ), .C2(n225), .ZN(n240) );
  AOI22_X2 U36 ( .A1(\U26/DATA1_4 ), .A2(n222), .B1(ElementAddr[4]), .B2(n223), 
        .ZN(n237) );
  AOI222_X1 U37 ( .A1(\U23/DATA1_4 ), .A2(n232), .B1(\U26/DATA2_4 ), .B2(n874), 
        .C1(\U20/DATA1_4 ), .C2(n225), .ZN(n238) );
  AOI22_X2 U38 ( .A1(\U26/DATA1_5 ), .A2(n222), .B1(ElementAddr[5]), .B2(n223), 
        .ZN(n235) );
  AOI222_X1 U39 ( .A1(\U23/DATA1_5 ), .A2(n232), .B1(\U26/DATA2_5 ), .B2(n874), 
        .C1(\U20/DATA1_5 ), .C2(n225), .ZN(n236) );
  AOI22_X2 U40 ( .A1(\U26/DATA1_6 ), .A2(n222), .B1(ElementAddr[6]), .B2(n223), 
        .ZN(n233) );
  AOI222_X1 U41 ( .A1(\U23/DATA1_6 ), .A2(n232), .B1(\U26/DATA2_6 ), .B2(n874), 
        .C1(\U20/DATA1_6 ), .C2(n225), .ZN(n234) );
  AOI22_X2 U42 ( .A1(\U26/DATA1_7 ), .A2(n222), .B1(ElementAddr[7]), .B2(n223), 
        .ZN(n230) );
  AOI222_X1 U43 ( .A1(\U23/DATA1_7 ), .A2(n232), .B1(\U26/DATA2_7 ), .B2(n874), 
        .C1(\U20/DATA1_7 ), .C2(n225), .ZN(n231) );
  OAI211_X2 U44 ( .C1(n869), .C2(n945), .A(n343), .B(n344), .ZN(n475) );
  AOI22_X2 U45 ( .A1(\U27/DATA1_47 ), .A2(n876), .B1(Element[47]), .B2(n866), 
        .ZN(n344) );
  AOI22_X2 U46 ( .A1(n874), .A2(\U27/DATA2_47 ), .B1(\U21/DATA1_47 ), .B2(n225), .ZN(n343) );
  OAI211_X2 U47 ( .C1(n870), .C2(n946), .A(n341), .B(n342), .ZN(n474) );
  AOI22_X2 U48 ( .A1(\U27/DATA1_46 ), .A2(n876), .B1(Element[46]), .B2(n866), 
        .ZN(n342) );
  AOI22_X2 U49 ( .A1(n874), .A2(\U27/DATA2_46 ), .B1(\U21/DATA1_46 ), .B2(n872), .ZN(n341) );
  OAI211_X2 U50 ( .C1(n869), .C2(n947), .A(n339), .B(n340), .ZN(n473) );
  AOI22_X2 U51 ( .A1(\U27/DATA1_45 ), .A2(n876), .B1(Element[45]), .B2(n866), 
        .ZN(n340) );
  AOI22_X2 U52 ( .A1(n874), .A2(\U27/DATA2_45 ), .B1(\U21/DATA1_45 ), .B2(n872), .ZN(n339) );
  OAI211_X2 U53 ( .C1(n870), .C2(n948), .A(n337), .B(n338), .ZN(n472) );
  AOI22_X2 U54 ( .A1(\U27/DATA1_44 ), .A2(n876), .B1(Element[44]), .B2(n866), 
        .ZN(n338) );
  AOI22_X2 U55 ( .A1(n224), .A2(\U27/DATA2_44 ), .B1(\U21/DATA1_44 ), .B2(n872), .ZN(n337) );
  OAI211_X2 U56 ( .C1(n869), .C2(n949), .A(n335), .B(n336), .ZN(n471) );
  AOI22_X2 U57 ( .A1(\U27/DATA1_43 ), .A2(n876), .B1(Element[43]), .B2(n866), 
        .ZN(n336) );
  AOI22_X2 U58 ( .A1(n224), .A2(\U27/DATA2_43 ), .B1(\U21/DATA1_43 ), .B2(n872), .ZN(n335) );
  OAI211_X2 U59 ( .C1(n870), .C2(n950), .A(n333), .B(n334), .ZN(n470) );
  AOI22_X2 U60 ( .A1(\U27/DATA1_42 ), .A2(n876), .B1(Element[42]), .B2(n866), 
        .ZN(n334) );
  AOI22_X2 U61 ( .A1(n874), .A2(\U27/DATA2_42 ), .B1(\U21/DATA1_42 ), .B2(n872), .ZN(n333) );
  OAI211_X2 U62 ( .C1(n869), .C2(n951), .A(n331), .B(n332), .ZN(n469) );
  AOI22_X2 U63 ( .A1(\U27/DATA1_41 ), .A2(n876), .B1(Element[41]), .B2(n866), 
        .ZN(n332) );
  AOI22_X2 U64 ( .A1(n224), .A2(\U27/DATA2_41 ), .B1(\U21/DATA1_41 ), .B2(n872), .ZN(n331) );
  OAI211_X2 U65 ( .C1(n869), .C2(n952), .A(n329), .B(n330), .ZN(n468) );
  AOI22_X2 U66 ( .A1(\U27/DATA1_40 ), .A2(n876), .B1(Element[40]), .B2(n866), 
        .ZN(n330) );
  AOI22_X2 U67 ( .A1(n874), .A2(\U27/DATA2_40 ), .B1(\U21/DATA1_40 ), .B2(n872), .ZN(n329) );
  OAI211_X2 U68 ( .C1(n870), .C2(n953), .A(n327), .B(n328), .ZN(n467) );
  AOI22_X2 U69 ( .A1(\U27/DATA1_39 ), .A2(n876), .B1(Element[39]), .B2(n866), 
        .ZN(n328) );
  AOI22_X2 U70 ( .A1(n224), .A2(\U27/DATA2_39 ), .B1(\U21/DATA1_39 ), .B2(n872), .ZN(n327) );
  OAI211_X2 U71 ( .C1(n870), .C2(n954), .A(n325), .B(n326), .ZN(n466) );
  AOI22_X2 U72 ( .A1(\U27/DATA1_38 ), .A2(n876), .B1(Element[38]), .B2(n866), 
        .ZN(n326) );
  AOI22_X2 U73 ( .A1(n874), .A2(\U27/DATA2_38 ), .B1(\U21/DATA1_38 ), .B2(n872), .ZN(n325) );
  OAI211_X2 U74 ( .C1(n869), .C2(n955), .A(n323), .B(n324), .ZN(n465) );
  AOI22_X2 U75 ( .A1(\U27/DATA1_37 ), .A2(n876), .B1(Element[37]), .B2(n866), 
        .ZN(n324) );
  AOI22_X2 U76 ( .A1(n224), .A2(\U27/DATA2_37 ), .B1(\U21/DATA1_37 ), .B2(n872), .ZN(n323) );
  OAI211_X2 U77 ( .C1(n870), .C2(n956), .A(n321), .B(n322), .ZN(n464) );
  AOI22_X2 U78 ( .A1(\U27/DATA1_36 ), .A2(n876), .B1(Element[36]), .B2(n866), 
        .ZN(n322) );
  AOI22_X2 U79 ( .A1(n874), .A2(\U27/DATA2_36 ), .B1(\U21/DATA1_36 ), .B2(n872), .ZN(n321) );
  OAI211_X2 U80 ( .C1(n869), .C2(n957), .A(n319), .B(n320), .ZN(n463) );
  AOI22_X2 U81 ( .A1(\U27/DATA1_35 ), .A2(n877), .B1(Element[35]), .B2(n866), 
        .ZN(n320) );
  AOI22_X2 U82 ( .A1(n224), .A2(\U27/DATA2_35 ), .B1(\U21/DATA1_35 ), .B2(n872), .ZN(n319) );
  OAI211_X2 U83 ( .C1(n869), .C2(n958), .A(n317), .B(n318), .ZN(n462) );
  AOI22_X2 U84 ( .A1(\U27/DATA1_34 ), .A2(n877), .B1(Element[34]), .B2(n866), 
        .ZN(n318) );
  AOI22_X2 U85 ( .A1(n874), .A2(\U27/DATA2_34 ), .B1(\U21/DATA1_34 ), .B2(n872), .ZN(n317) );
  OAI211_X2 U86 ( .C1(n869), .C2(n959), .A(n315), .B(n316), .ZN(n461) );
  AOI22_X2 U87 ( .A1(\U27/DATA1_33 ), .A2(n877), .B1(Element[33]), .B2(n866), 
        .ZN(n316) );
  AOI22_X2 U88 ( .A1(n224), .A2(\U27/DATA2_33 ), .B1(\U21/DATA1_33 ), .B2(n872), .ZN(n315) );
  OAI211_X2 U89 ( .C1(n869), .C2(n960), .A(n313), .B(n314), .ZN(n460) );
  AOI22_X2 U90 ( .A1(\U27/DATA1_32 ), .A2(n877), .B1(Element[32]), .B2(n866), 
        .ZN(n314) );
  AOI22_X2 U91 ( .A1(n874), .A2(\U27/DATA2_32 ), .B1(\U21/DATA1_32 ), .B2(n872), .ZN(n313) );
  OAI211_X2 U92 ( .C1(n869), .C2(n961), .A(n311), .B(n312), .ZN(n459) );
  AOI22_X2 U93 ( .A1(\U27/DATA1_31 ), .A2(n877), .B1(Element[31]), .B2(n866), 
        .ZN(n312) );
  AOI22_X2 U94 ( .A1(n874), .A2(\U27/DATA2_31 ), .B1(\U21/DATA1_31 ), .B2(n872), .ZN(n311) );
  OAI211_X2 U95 ( .C1(n869), .C2(n962), .A(n309), .B(n310), .ZN(n458) );
  AOI22_X2 U96 ( .A1(\U27/DATA1_30 ), .A2(n877), .B1(Element[30]), .B2(n866), 
        .ZN(n310) );
  AOI22_X2 U97 ( .A1(n874), .A2(\U27/DATA2_30 ), .B1(\U21/DATA1_30 ), .B2(n872), .ZN(n309) );
  OAI211_X2 U98 ( .C1(n869), .C2(n963), .A(n307), .B(n308), .ZN(n457) );
  AOI22_X2 U99 ( .A1(\U27/DATA1_29 ), .A2(n877), .B1(Element[29]), .B2(n866), 
        .ZN(n308) );
  AOI22_X2 U100 ( .A1(n874), .A2(\U27/DATA2_29 ), .B1(\U21/DATA1_29 ), .B2(
        n872), .ZN(n307) );
  OAI211_X2 U101 ( .C1(n869), .C2(n964), .A(n305), .B(n306), .ZN(n456) );
  AOI22_X2 U102 ( .A1(\U27/DATA1_28 ), .A2(n877), .B1(Element[28]), .B2(n866), 
        .ZN(n306) );
  AOI22_X2 U103 ( .A1(n874), .A2(\U27/DATA2_28 ), .B1(\U21/DATA1_28 ), .B2(
        n225), .ZN(n305) );
  OAI211_X2 U104 ( .C1(n869), .C2(n965), .A(n303), .B(n304), .ZN(n455) );
  AOI22_X2 U105 ( .A1(\U27/DATA1_27 ), .A2(n877), .B1(Element[27]), .B2(n866), 
        .ZN(n304) );
  AOI22_X2 U106 ( .A1(n874), .A2(\U27/DATA2_27 ), .B1(\U21/DATA1_27 ), .B2(
        n225), .ZN(n303) );
  OAI211_X2 U107 ( .C1(n869), .C2(n966), .A(n301), .B(n302), .ZN(n454) );
  AOI22_X2 U108 ( .A1(\U27/DATA1_26 ), .A2(n877), .B1(Element[26]), .B2(n866), 
        .ZN(n302) );
  AOI22_X2 U109 ( .A1(n874), .A2(\U27/DATA2_26 ), .B1(\U21/DATA1_26 ), .B2(
        n225), .ZN(n301) );
  OAI211_X2 U110 ( .C1(n869), .C2(n967), .A(n299), .B(n300), .ZN(n453) );
  AOI22_X2 U111 ( .A1(\U27/DATA1_25 ), .A2(n877), .B1(Element[25]), .B2(n866), 
        .ZN(n300) );
  AOI22_X2 U112 ( .A1(n874), .A2(\U27/DATA2_25 ), .B1(\U21/DATA1_25 ), .B2(
        n225), .ZN(n299) );
  OAI211_X2 U113 ( .C1(n869), .C2(n968), .A(n297), .B(n298), .ZN(n452) );
  AOI22_X2 U114 ( .A1(\U27/DATA1_24 ), .A2(n877), .B1(Element[24]), .B2(n866), 
        .ZN(n298) );
  AOI22_X2 U115 ( .A1(n874), .A2(\U27/DATA2_24 ), .B1(\U21/DATA1_24 ), .B2(
        n225), .ZN(n297) );
  OAI211_X2 U116 ( .C1(n869), .C2(n969), .A(n295), .B(n296), .ZN(n451) );
  AOI22_X2 U117 ( .A1(\U27/DATA1_23 ), .A2(n876), .B1(Element[23]), .B2(n866), 
        .ZN(n296) );
  AOI22_X2 U118 ( .A1(n874), .A2(\U27/DATA2_23 ), .B1(\U21/DATA1_23 ), .B2(
        n225), .ZN(n295) );
  OAI211_X2 U119 ( .C1(n869), .C2(n970), .A(n293), .B(n294), .ZN(n450) );
  AOI22_X2 U120 ( .A1(\U27/DATA1_22 ), .A2(n877), .B1(Element[22]), .B2(n866), 
        .ZN(n294) );
  AOI22_X2 U121 ( .A1(n874), .A2(\U27/DATA2_22 ), .B1(\U21/DATA1_22 ), .B2(
        n225), .ZN(n293) );
  OAI211_X2 U122 ( .C1(n870), .C2(n971), .A(n291), .B(n292), .ZN(n449) );
  AOI22_X2 U123 ( .A1(\U27/DATA1_21 ), .A2(n222), .B1(Element[21]), .B2(n866), 
        .ZN(n292) );
  AOI22_X2 U124 ( .A1(n874), .A2(\U27/DATA2_21 ), .B1(\U21/DATA1_21 ), .B2(
        n225), .ZN(n291) );
  OAI211_X2 U125 ( .C1(n870), .C2(n972), .A(n289), .B(n290), .ZN(n448) );
  AOI22_X2 U126 ( .A1(\U27/DATA1_20 ), .A2(n222), .B1(Element[20]), .B2(n866), 
        .ZN(n290) );
  AOI22_X2 U127 ( .A1(n874), .A2(\U27/DATA2_20 ), .B1(\U21/DATA1_20 ), .B2(
        n225), .ZN(n289) );
  OAI211_X2 U128 ( .C1(n870), .C2(n973), .A(n287), .B(n288), .ZN(n447) );
  AOI22_X2 U129 ( .A1(\U27/DATA1_19 ), .A2(n222), .B1(Element[19]), .B2(n866), 
        .ZN(n288) );
  AOI22_X2 U130 ( .A1(n874), .A2(\U27/DATA2_19 ), .B1(\U21/DATA1_19 ), .B2(
        n225), .ZN(n287) );
  OAI211_X2 U131 ( .C1(n870), .C2(n974), .A(n285), .B(n286), .ZN(n446) );
  AOI22_X2 U132 ( .A1(\U27/DATA1_18 ), .A2(n222), .B1(Element[18]), .B2(n866), 
        .ZN(n286) );
  AOI22_X2 U133 ( .A1(n874), .A2(\U27/DATA2_18 ), .B1(\U21/DATA1_18 ), .B2(
        n225), .ZN(n285) );
  OAI211_X2 U134 ( .C1(n870), .C2(n975), .A(n283), .B(n284), .ZN(n445) );
  AOI22_X2 U135 ( .A1(\U27/DATA1_17 ), .A2(n222), .B1(Element[17]), .B2(n866), 
        .ZN(n284) );
  AOI22_X2 U136 ( .A1(n874), .A2(\U27/DATA2_17 ), .B1(\U21/DATA1_17 ), .B2(
        n225), .ZN(n283) );
  OAI211_X2 U137 ( .C1(n870), .C2(n976), .A(n281), .B(n282), .ZN(n444) );
  AOI22_X2 U138 ( .A1(\U27/DATA1_16 ), .A2(n222), .B1(Element[16]), .B2(n866), 
        .ZN(n282) );
  AOI22_X2 U139 ( .A1(n224), .A2(\U27/DATA2_16 ), .B1(\U21/DATA1_16 ), .B2(
        n872), .ZN(n281) );
  OAI211_X2 U140 ( .C1(n870), .C2(n977), .A(n279), .B(n280), .ZN(n443) );
  AOI22_X2 U141 ( .A1(\U27/DATA1_15 ), .A2(n222), .B1(Element[15]), .B2(n866), 
        .ZN(n280) );
  AOI22_X2 U142 ( .A1(n224), .A2(\U27/DATA2_15 ), .B1(\U21/DATA1_15 ), .B2(
        n872), .ZN(n279) );
  OAI211_X2 U143 ( .C1(n870), .C2(n978), .A(n277), .B(n278), .ZN(n442) );
  AOI22_X2 U144 ( .A1(\U27/DATA1_14 ), .A2(n222), .B1(Element[14]), .B2(n866), 
        .ZN(n278) );
  AOI22_X2 U145 ( .A1(n224), .A2(\U27/DATA2_14 ), .B1(\U21/DATA1_14 ), .B2(
        n872), .ZN(n277) );
  OAI211_X2 U146 ( .C1(n870), .C2(n979), .A(n275), .B(n276), .ZN(n441) );
  AOI22_X2 U147 ( .A1(\U27/DATA1_13 ), .A2(n222), .B1(Element[13]), .B2(n866), 
        .ZN(n276) );
  AOI22_X2 U148 ( .A1(n224), .A2(\U27/DATA2_13 ), .B1(\U21/DATA1_13 ), .B2(
        n872), .ZN(n275) );
  OAI211_X2 U149 ( .C1(n870), .C2(n980), .A(n273), .B(n274), .ZN(n440) );
  AOI22_X2 U150 ( .A1(\U27/DATA1_12 ), .A2(n222), .B1(Element[12]), .B2(n866), 
        .ZN(n274) );
  AOI22_X2 U151 ( .A1(n224), .A2(\U27/DATA2_12 ), .B1(\U21/DATA1_12 ), .B2(
        n225), .ZN(n273) );
  OAI211_X2 U152 ( .C1(n870), .C2(n981), .A(n271), .B(n272), .ZN(n439) );
  AOI22_X2 U153 ( .A1(\U27/DATA1_11 ), .A2(n876), .B1(Element[11]), .B2(n866), 
        .ZN(n272) );
  AOI22_X2 U154 ( .A1(n224), .A2(\U27/DATA2_11 ), .B1(\U21/DATA1_11 ), .B2(
        n872), .ZN(n271) );
  OAI211_X2 U155 ( .C1(n870), .C2(n982), .A(n269), .B(n270), .ZN(n438) );
  AOI22_X2 U157 ( .A1(\U27/DATA1_10 ), .A2(n876), .B1(Element[10]), .B2(n866), 
        .ZN(n270) );
  AOI22_X2 U158 ( .A1(n224), .A2(\U27/DATA2_10 ), .B1(\U21/DATA1_10 ), .B2(
        n872), .ZN(n269) );
  OAI211_X2 U160 ( .C1(n870), .C2(n983), .A(n267), .B(n268), .ZN(n437) );
  AOI22_X2 U161 ( .A1(\U27/DATA1_9 ), .A2(n877), .B1(Element[9]), .B2(n866), 
        .ZN(n268) );
  AOI22_X2 U163 ( .A1(n224), .A2(\U27/DATA2_9 ), .B1(\U21/DATA1_9 ), .B2(n872), 
        .ZN(n267) );
  OAI211_X2 U164 ( .C1(n869), .C2(n984), .A(n265), .B(n266), .ZN(n436) );
  AOI22_X2 U166 ( .A1(\U27/DATA1_8 ), .A2(n877), .B1(Element[8]), .B2(n866), 
        .ZN(n266) );
  AOI22_X2 U167 ( .A1(n224), .A2(\U27/DATA2_8 ), .B1(\U21/DATA1_8 ), .B2(n872), 
        .ZN(n265) );
  OAI211_X2 U169 ( .C1(n870), .C2(n985), .A(n263), .B(n264), .ZN(n435) );
  AOI22_X2 U170 ( .A1(\U27/DATA1_7 ), .A2(n876), .B1(Element[7]), .B2(n866), 
        .ZN(n264) );
  AOI22_X2 U172 ( .A1(n224), .A2(\U27/DATA2_7 ), .B1(\U21/DATA1_7 ), .B2(n872), 
        .ZN(n263) );
  OAI211_X2 U173 ( .C1(n870), .C2(n986), .A(n261), .B(n262), .ZN(n434) );
  AOI22_X2 U175 ( .A1(\U27/DATA1_6 ), .A2(n877), .B1(Element[6]), .B2(n866), 
        .ZN(n262) );
  AOI22_X2 U176 ( .A1(n224), .A2(\U27/DATA2_6 ), .B1(\U21/DATA1_6 ), .B2(n872), 
        .ZN(n261) );
  OAI211_X2 U178 ( .C1(n869), .C2(n987), .A(n259), .B(n260), .ZN(n433) );
  AOI22_X2 U179 ( .A1(\U27/DATA1_5 ), .A2(n222), .B1(Element[5]), .B2(n866), 
        .ZN(n260) );
  AOI22_X2 U180 ( .A1(n224), .A2(\U27/DATA2_5 ), .B1(\U21/DATA1_5 ), .B2(n872), 
        .ZN(n259) );
  OAI211_X2 U181 ( .C1(n870), .C2(n988), .A(n257), .B(n258), .ZN(n432) );
  AOI22_X2 U182 ( .A1(\U27/DATA1_4 ), .A2(n222), .B1(Element[4]), .B2(n866), 
        .ZN(n258) );
  AOI22_X2 U183 ( .A1(n874), .A2(\U27/DATA2_4 ), .B1(\U21/DATA1_4 ), .B2(n872), 
        .ZN(n257) );
  OAI211_X2 U184 ( .C1(n869), .C2(n989), .A(n255), .B(n256), .ZN(n431) );
  AOI22_X2 U185 ( .A1(\U27/DATA1_3 ), .A2(n222), .B1(Element[3]), .B2(n866), 
        .ZN(n256) );
  AOI22_X2 U186 ( .A1(n874), .A2(\U27/DATA2_3 ), .B1(\U21/DATA1_3 ), .B2(n225), 
        .ZN(n255) );
  OAI211_X2 U187 ( .C1(n870), .C2(n990), .A(n253), .B(n254), .ZN(n430) );
  AOI22_X2 U188 ( .A1(\U27/DATA1_2 ), .A2(n222), .B1(Element[2]), .B2(n866), 
        .ZN(n254) );
  AOI22_X2 U189 ( .A1(n874), .A2(\U27/DATA2_2 ), .B1(\U21/DATA1_2 ), .B2(n225), 
        .ZN(n253) );
  OAI211_X2 U190 ( .C1(n869), .C2(n991), .A(n251), .B(n252), .ZN(n429) );
  AOI22_X2 U191 ( .A1(\U27/DATA1_1 ), .A2(n222), .B1(Element[1]), .B2(n866), 
        .ZN(n252) );
  AOI22_X2 U192 ( .A1(n874), .A2(\U27/DATA2_1 ), .B1(\U21/DATA1_1 ), .B2(n225), 
        .ZN(n251) );
  OAI211_X2 U193 ( .C1(n870), .C2(n992), .A(n248), .B(n249), .ZN(n428) );
  AOI22_X2 U194 ( .A1(\U27/DATA1_0 ), .A2(n222), .B1(Element[0]), .B2(n866), 
        .ZN(n249) );
  AOI22_X2 U195 ( .A1(n874), .A2(\U27/DATA2_0 ), .B1(\U21/DATA1_0 ), .B2(n872), 
        .ZN(n248) );
  OAI211_X2 U196 ( .C1(n869), .C2(n944), .A(n228), .B(n229), .ZN(n419) );
  AOI22_X2 U197 ( .A1(\U3/U5/DATA2_0 ), .A2(n876), .B1(ElementAddr[8]), .B2(
        n223), .ZN(n229) );
  AOI22_X2 U198 ( .A1(\U3/U5/DATA3_0 ), .A2(n874), .B1(\U20/DATA1_8 ), .B2(
        n225), .ZN(n228) );
  OAI211_X2 U199 ( .C1(n870), .C2(n943), .A(n226), .B(n227), .ZN(n418) );
  AOI22_X2 U200 ( .A1(\U3/U5/DATA2_1 ), .A2(n877), .B1(ElementAddr[9]), .B2(
        n223), .ZN(n227) );
  AOI22_X2 U201 ( .A1(\U3/U5/DATA3_1 ), .A2(n874), .B1(\U20/DATA1_9 ), .B2(
        n872), .ZN(n226) );
  OAI211_X2 U202 ( .C1(n869), .C2(n942), .A(n220), .B(n221), .ZN(n417) );
  AOI22_X2 U203 ( .A1(\U3/U5/DATA2_2 ), .A2(n222), .B1(ElementAddr[10]), .B2(
        n223), .ZN(n221) );
  AOI22_X2 U204 ( .A1(\U3/U5/DATA3_2 ), .A2(n874), .B1(\U20/DATA1_10 ), .B2(
        n225), .ZN(n220) );
  OAI222_X2 U205 ( .A1(n247), .A2(n358), .B1(n359), .B2(n891), .C1(n868), .C2(
        n994), .ZN(n480) );
  AOI21_X2 U206 ( .B1(\r389/A[2] ), .B2(n893), .A(n360), .ZN(n359) );
  OAI222_X2 U207 ( .A1(n354), .A2(n891), .B1(n355), .B2(n247), .C1(n868), .C2(
        n995), .ZN(n479) );
  AOI21_X2 U208 ( .B1(\r389/A[1] ), .B2(\r389/A[0] ), .A(n357), .ZN(n354) );
  AOI21_X2 U209 ( .B1(n884), .B2(n883), .A(n356), .ZN(n355) );
  OAI222_X2 U210 ( .A1(n868), .A2(n996), .B1(n883), .B2(n247), .C1(\r389/A[0] ), .C2(n891), .ZN(n478) );
  OAI211_X2 U211 ( .C1(n120), .C2(n918), .A(n171), .B(n172), .ZN(n393) );
  AOI22_X2 U212 ( .A1(\U27/DATA2_23 ), .A2(n871), .B1(\U24/DATA1_23 ), .B2(
        n879), .ZN(n171) );
  AOI22_X2 U213 ( .A1(\U21/DATA1_23 ), .A2(n880), .B1(Diagonal[23]), .B2(n888), 
        .ZN(n172) );
  OAI211_X2 U214 ( .C1(n120), .C2(n905), .A(n145), .B(n146), .ZN(n380) );
  AOI22_X2 U215 ( .A1(\U27/DATA2_36 ), .A2(n871), .B1(\U24/DATA1_36 ), .B2(
        n879), .ZN(n145) );
  AOI22_X2 U216 ( .A1(\U21/DATA1_36 ), .A2(n880), .B1(Diagonal[36]), .B2(n888), 
        .ZN(n146) );
  OAI211_X2 U217 ( .C1(n882), .C2(n904), .A(n143), .B(n144), .ZN(n379) );
  AOI22_X2 U218 ( .A1(\U27/DATA2_37 ), .A2(n871), .B1(\U24/DATA1_37 ), .B2(
        n879), .ZN(n143) );
  AOI22_X2 U219 ( .A1(\U21/DATA1_37 ), .A2(n880), .B1(Diagonal[37]), .B2(n888), 
        .ZN(n144) );
  OAI211_X2 U220 ( .C1(n120), .C2(n903), .A(n141), .B(n142), .ZN(n378) );
  AOI22_X2 U221 ( .A1(\U27/DATA2_38 ), .A2(n871), .B1(\U24/DATA1_38 ), .B2(
        n879), .ZN(n141) );
  AOI22_X2 U222 ( .A1(\U21/DATA1_38 ), .A2(n880), .B1(Diagonal[38]), .B2(n888), 
        .ZN(n142) );
  OAI211_X2 U223 ( .C1(n882), .C2(n902), .A(n139), .B(n140), .ZN(n377) );
  AOI22_X2 U224 ( .A1(\U27/DATA2_39 ), .A2(n871), .B1(\U24/DATA1_39 ), .B2(
        n879), .ZN(n139) );
  AOI22_X2 U225 ( .A1(\U21/DATA1_39 ), .A2(n880), .B1(Diagonal[39]), .B2(n888), 
        .ZN(n140) );
  OAI211_X2 U226 ( .C1(n120), .C2(n901), .A(n137), .B(n138), .ZN(n376) );
  AOI22_X2 U227 ( .A1(\U27/DATA2_40 ), .A2(n871), .B1(\U24/DATA1_40 ), .B2(
        n879), .ZN(n137) );
  AOI22_X2 U228 ( .A1(\U21/DATA1_40 ), .A2(n880), .B1(Diagonal[40]), .B2(n888), 
        .ZN(n138) );
  OAI211_X2 U229 ( .C1(n882), .C2(n900), .A(n135), .B(n136), .ZN(n375) );
  AOI22_X2 U230 ( .A1(\U27/DATA2_41 ), .A2(n871), .B1(\U24/DATA1_41 ), .B2(
        n879), .ZN(n135) );
  AOI22_X2 U231 ( .A1(\U21/DATA1_41 ), .A2(n880), .B1(Diagonal[41]), .B2(n888), 
        .ZN(n136) );
  OAI211_X2 U232 ( .C1(n120), .C2(n899), .A(n133), .B(n134), .ZN(n374) );
  AOI22_X2 U233 ( .A1(\U27/DATA2_42 ), .A2(n871), .B1(\U24/DATA1_42 ), .B2(
        n879), .ZN(n133) );
  AOI22_X2 U234 ( .A1(\U21/DATA1_42 ), .A2(n880), .B1(Diagonal[42]), .B2(n888), 
        .ZN(n134) );
  OAI211_X2 U235 ( .C1(n120), .C2(n898), .A(n131), .B(n132), .ZN(n373) );
  AOI22_X2 U236 ( .A1(\U27/DATA2_43 ), .A2(n871), .B1(\U24/DATA1_43 ), .B2(
        n879), .ZN(n131) );
  AOI22_X2 U237 ( .A1(\U21/DATA1_43 ), .A2(n880), .B1(Diagonal[43]), .B2(n888), 
        .ZN(n132) );
  OAI211_X2 U238 ( .C1(n120), .C2(n897), .A(n129), .B(n130), .ZN(n372) );
  AOI22_X2 U239 ( .A1(\U27/DATA2_44 ), .A2(n871), .B1(\U24/DATA1_44 ), .B2(
        n879), .ZN(n129) );
  AOI22_X2 U240 ( .A1(\U21/DATA1_44 ), .A2(n880), .B1(Diagonal[44]), .B2(n888), 
        .ZN(n130) );
  OAI211_X2 U241 ( .C1(n120), .C2(n896), .A(n127), .B(n128), .ZN(n371) );
  AOI22_X2 U242 ( .A1(\U27/DATA2_45 ), .A2(n871), .B1(\U24/DATA1_45 ), .B2(
        n879), .ZN(n127) );
  AOI22_X2 U243 ( .A1(\U21/DATA1_45 ), .A2(n880), .B1(Diagonal[45]), .B2(n888), 
        .ZN(n128) );
  OAI211_X2 U244 ( .C1(n120), .C2(n895), .A(n125), .B(n126), .ZN(n370) );
  AOI22_X2 U245 ( .A1(\U27/DATA2_46 ), .A2(n871), .B1(\U24/DATA1_46 ), .B2(
        n879), .ZN(n125) );
  AOI22_X2 U246 ( .A1(\U21/DATA1_46 ), .A2(n880), .B1(Diagonal[46]), .B2(n888), 
        .ZN(n126) );
  OAI211_X2 U247 ( .C1(n882), .C2(n941), .A(n217), .B(n218), .ZN(n416) );
  AOI22_X2 U248 ( .A1(\U27/DATA2_0 ), .A2(n871), .B1(\U24/DATA1_0 ), .B2(n879), 
        .ZN(n217) );
  AOI22_X2 U249 ( .A1(\U21/DATA1_0 ), .A2(n880), .B1(Diagonal[0]), .B2(n888), 
        .ZN(n218) );
  OAI211_X2 U250 ( .C1(n882), .C2(n940), .A(n215), .B(n216), .ZN(n415) );
  AOI22_X2 U251 ( .A1(\U27/DATA2_1 ), .A2(n871), .B1(\U24/DATA1_1 ), .B2(n879), 
        .ZN(n215) );
  AOI22_X2 U252 ( .A1(\U21/DATA1_1 ), .A2(n880), .B1(Diagonal[1]), .B2(n888), 
        .ZN(n216) );
  OAI211_X2 U253 ( .C1(n882), .C2(n939), .A(n213), .B(n214), .ZN(n414) );
  AOI22_X2 U254 ( .A1(\U27/DATA2_2 ), .A2(n871), .B1(\U24/DATA1_2 ), .B2(n879), 
        .ZN(n213) );
  AOI22_X2 U255 ( .A1(\U21/DATA1_2 ), .A2(n880), .B1(Diagonal[2]), .B2(n888), 
        .ZN(n214) );
  OAI211_X2 U256 ( .C1(n882), .C2(n938), .A(n211), .B(n212), .ZN(n413) );
  AOI22_X2 U257 ( .A1(\U27/DATA2_3 ), .A2(n871), .B1(\U24/DATA1_3 ), .B2(n879), 
        .ZN(n211) );
  AOI22_X2 U258 ( .A1(\U21/DATA1_3 ), .A2(n880), .B1(Diagonal[3]), .B2(n888), 
        .ZN(n212) );
  OAI211_X2 U259 ( .C1(n882), .C2(n937), .A(n209), .B(n210), .ZN(n412) );
  AOI22_X2 U260 ( .A1(\U27/DATA2_4 ), .A2(n871), .B1(\U24/DATA1_4 ), .B2(n879), 
        .ZN(n209) );
  AOI22_X2 U261 ( .A1(\U21/DATA1_4 ), .A2(n880), .B1(Diagonal[4]), .B2(n888), 
        .ZN(n210) );
  OAI211_X2 U262 ( .C1(n882), .C2(n936), .A(n207), .B(n208), .ZN(n411) );
  AOI22_X2 U263 ( .A1(\U27/DATA2_5 ), .A2(n871), .B1(\U24/DATA1_5 ), .B2(n879), 
        .ZN(n207) );
  AOI22_X2 U264 ( .A1(\U21/DATA1_5 ), .A2(n880), .B1(Diagonal[5]), .B2(n888), 
        .ZN(n208) );
  OAI211_X2 U265 ( .C1(n882), .C2(n935), .A(n205), .B(n206), .ZN(n410) );
  AOI22_X2 U266 ( .A1(\U27/DATA2_6 ), .A2(n871), .B1(\U24/DATA1_6 ), .B2(n879), 
        .ZN(n205) );
  AOI22_X2 U267 ( .A1(\U21/DATA1_6 ), .A2(n880), .B1(Diagonal[6]), .B2(n888), 
        .ZN(n206) );
  OAI211_X2 U268 ( .C1(n882), .C2(n934), .A(n203), .B(n204), .ZN(n409) );
  AOI22_X2 U269 ( .A1(\U27/DATA2_7 ), .A2(n871), .B1(\U24/DATA1_7 ), .B2(n879), 
        .ZN(n203) );
  AOI22_X2 U270 ( .A1(\U21/DATA1_7 ), .A2(n880), .B1(Diagonal[7]), .B2(n888), 
        .ZN(n204) );
  OAI211_X2 U271 ( .C1(n882), .C2(n933), .A(n201), .B(n202), .ZN(n408) );
  AOI22_X2 U272 ( .A1(\U27/DATA2_8 ), .A2(n871), .B1(\U24/DATA1_8 ), .B2(n879), 
        .ZN(n201) );
  AOI22_X2 U273 ( .A1(\U21/DATA1_8 ), .A2(n880), .B1(Diagonal[8]), .B2(n888), 
        .ZN(n202) );
  OAI211_X2 U274 ( .C1(n882), .C2(n932), .A(n199), .B(n200), .ZN(n407) );
  AOI22_X2 U275 ( .A1(\U27/DATA2_9 ), .A2(n871), .B1(\U24/DATA1_9 ), .B2(n879), 
        .ZN(n199) );
  AOI22_X2 U276 ( .A1(\U21/DATA1_9 ), .A2(n880), .B1(Diagonal[9]), .B2(n888), 
        .ZN(n200) );
  OAI211_X2 U277 ( .C1(n882), .C2(n931), .A(n197), .B(n198), .ZN(n406) );
  AOI22_X2 U278 ( .A1(\U27/DATA2_10 ), .A2(n871), .B1(\U24/DATA1_10 ), .B2(
        n879), .ZN(n197) );
  AOI22_X2 U279 ( .A1(\U21/DATA1_10 ), .A2(n880), .B1(Diagonal[10]), .B2(n888), 
        .ZN(n198) );
  OAI211_X2 U280 ( .C1(n882), .C2(n930), .A(n195), .B(n196), .ZN(n405) );
  AOI22_X2 U281 ( .A1(\U27/DATA2_11 ), .A2(n871), .B1(\U24/DATA1_11 ), .B2(
        n879), .ZN(n195) );
  AOI22_X2 U282 ( .A1(\U21/DATA1_11 ), .A2(n880), .B1(Diagonal[11]), .B2(n888), 
        .ZN(n196) );
  OAI211_X2 U283 ( .C1(n882), .C2(n929), .A(n193), .B(n194), .ZN(n404) );
  AOI22_X2 U284 ( .A1(\U27/DATA2_12 ), .A2(n871), .B1(\U24/DATA1_12 ), .B2(
        n879), .ZN(n193) );
  AOI22_X2 U285 ( .A1(\U21/DATA1_12 ), .A2(n880), .B1(Diagonal[12]), .B2(n888), 
        .ZN(n194) );
  OAI211_X2 U286 ( .C1(n882), .C2(n928), .A(n191), .B(n192), .ZN(n403) );
  AOI22_X2 U287 ( .A1(\U27/DATA2_13 ), .A2(n871), .B1(\U24/DATA1_13 ), .B2(
        n879), .ZN(n191) );
  AOI22_X2 U288 ( .A1(\U21/DATA1_13 ), .A2(n880), .B1(Diagonal[13]), .B2(n888), 
        .ZN(n192) );
  OAI211_X2 U289 ( .C1(n882), .C2(n927), .A(n189), .B(n190), .ZN(n402) );
  AOI22_X2 U290 ( .A1(\U27/DATA2_14 ), .A2(n871), .B1(\U24/DATA1_14 ), .B2(
        n879), .ZN(n189) );
  AOI22_X2 U291 ( .A1(\U21/DATA1_14 ), .A2(n880), .B1(Diagonal[14]), .B2(n888), 
        .ZN(n190) );
  OAI211_X2 U292 ( .C1(n882), .C2(n926), .A(n187), .B(n188), .ZN(n401) );
  AOI22_X2 U293 ( .A1(\U27/DATA2_15 ), .A2(n871), .B1(\U24/DATA1_15 ), .B2(
        n879), .ZN(n187) );
  AOI22_X2 U294 ( .A1(\U21/DATA1_15 ), .A2(n880), .B1(Diagonal[15]), .B2(n888), 
        .ZN(n188) );
  OAI211_X2 U295 ( .C1(n882), .C2(n925), .A(n185), .B(n186), .ZN(n400) );
  AOI22_X2 U296 ( .A1(\U27/DATA2_16 ), .A2(n871), .B1(\U24/DATA1_16 ), .B2(
        n879), .ZN(n185) );
  AOI22_X2 U297 ( .A1(\U21/DATA1_16 ), .A2(n880), .B1(Diagonal[16]), .B2(n888), 
        .ZN(n186) );
  OAI211_X2 U298 ( .C1(n882), .C2(n924), .A(n183), .B(n184), .ZN(n399) );
  AOI22_X2 U299 ( .A1(\U27/DATA2_17 ), .A2(n871), .B1(\U24/DATA1_17 ), .B2(
        n879), .ZN(n183) );
  AOI22_X2 U300 ( .A1(\U21/DATA1_17 ), .A2(n880), .B1(Diagonal[17]), .B2(n888), 
        .ZN(n184) );
  OAI211_X2 U301 ( .C1(n882), .C2(n923), .A(n181), .B(n182), .ZN(n398) );
  AOI22_X2 U302 ( .A1(\U27/DATA2_18 ), .A2(n871), .B1(\U24/DATA1_18 ), .B2(
        n879), .ZN(n181) );
  AOI22_X2 U303 ( .A1(\U21/DATA1_18 ), .A2(n880), .B1(Diagonal[18]), .B2(n888), 
        .ZN(n182) );
  OAI211_X2 U304 ( .C1(n882), .C2(n922), .A(n179), .B(n180), .ZN(n397) );
  AOI22_X2 U305 ( .A1(\U27/DATA2_19 ), .A2(n871), .B1(\U24/DATA1_19 ), .B2(
        n879), .ZN(n179) );
  AOI22_X2 U306 ( .A1(\U21/DATA1_19 ), .A2(n880), .B1(Diagonal[19]), .B2(n888), 
        .ZN(n180) );
  OAI211_X2 U307 ( .C1(n882), .C2(n921), .A(n177), .B(n178), .ZN(n396) );
  AOI22_X2 U308 ( .A1(\U27/DATA2_20 ), .A2(n871), .B1(\U24/DATA1_20 ), .B2(
        n879), .ZN(n177) );
  AOI22_X2 U309 ( .A1(\U21/DATA1_20 ), .A2(n880), .B1(Diagonal[20]), .B2(n888), 
        .ZN(n178) );
  OAI211_X2 U310 ( .C1(n882), .C2(n920), .A(n175), .B(n176), .ZN(n395) );
  AOI22_X2 U311 ( .A1(\U27/DATA2_21 ), .A2(n871), .B1(\U24/DATA1_21 ), .B2(
        n879), .ZN(n175) );
  AOI22_X2 U312 ( .A1(\U21/DATA1_21 ), .A2(n880), .B1(Diagonal[21]), .B2(n888), 
        .ZN(n176) );
  OAI211_X2 U313 ( .C1(n120), .C2(n919), .A(n173), .B(n174), .ZN(n394) );
  AOI22_X2 U314 ( .A1(\U27/DATA2_22 ), .A2(n871), .B1(\U24/DATA1_22 ), .B2(
        n879), .ZN(n173) );
  AOI22_X2 U315 ( .A1(\U21/DATA1_22 ), .A2(n880), .B1(Diagonal[22]), .B2(n888), 
        .ZN(n174) );
  OAI211_X2 U316 ( .C1(n120), .C2(n894), .A(n121), .B(n122), .ZN(n369) );
  AOI22_X2 U317 ( .A1(\U27/DATA2_47 ), .A2(n871), .B1(\U24/DATA1_47 ), .B2(
        n879), .ZN(n121) );
  AOI22_X2 U318 ( .A1(\U21/DATA1_47 ), .A2(n880), .B1(Diagonal[47]), .B2(n888), 
        .ZN(n122) );
  OAI211_X2 U319 ( .C1(n120), .C2(n917), .A(n169), .B(n170), .ZN(n392) );
  AOI22_X2 U320 ( .A1(\U27/DATA2_24 ), .A2(n871), .B1(\U24/DATA1_24 ), .B2(
        n879), .ZN(n169) );
  AOI22_X2 U321 ( .A1(\U21/DATA1_24 ), .A2(n880), .B1(Diagonal[24]), .B2(n888), 
        .ZN(n170) );
  OAI211_X2 U322 ( .C1(n120), .C2(n916), .A(n167), .B(n168), .ZN(n391) );
  AOI22_X2 U323 ( .A1(\U27/DATA2_25 ), .A2(n871), .B1(\U24/DATA1_25 ), .B2(
        n879), .ZN(n167) );
  AOI22_X2 U325 ( .A1(\U21/DATA1_25 ), .A2(n880), .B1(Diagonal[25]), .B2(n888), 
        .ZN(n168) );
  OAI211_X2 U326 ( .C1(n120), .C2(n915), .A(n165), .B(n166), .ZN(n390) );
  AOI22_X2 U327 ( .A1(\U27/DATA2_26 ), .A2(n871), .B1(\U24/DATA1_26 ), .B2(
        n879), .ZN(n165) );
  AOI22_X2 U329 ( .A1(\U21/DATA1_26 ), .A2(n880), .B1(Diagonal[26]), .B2(n888), 
        .ZN(n166) );
  OAI211_X2 U331 ( .C1(n120), .C2(n914), .A(n163), .B(n164), .ZN(n389) );
  AOI22_X2 U332 ( .A1(\U27/DATA2_27 ), .A2(n871), .B1(\U24/DATA1_27 ), .B2(
        n879), .ZN(n163) );
  AOI22_X2 U334 ( .A1(\U21/DATA1_27 ), .A2(n880), .B1(Diagonal[27]), .B2(n888), 
        .ZN(n164) );
  OAI211_X2 U336 ( .C1(n120), .C2(n913), .A(n161), .B(n162), .ZN(n388) );
  AOI22_X2 U337 ( .A1(\U27/DATA2_28 ), .A2(n871), .B1(\U24/DATA1_28 ), .B2(
        n879), .ZN(n161) );
  AOI22_X2 U338 ( .A1(\U21/DATA1_28 ), .A2(n880), .B1(Diagonal[28]), .B2(n888), 
        .ZN(n162) );
  OAI211_X2 U339 ( .C1(n120), .C2(n912), .A(n159), .B(n160), .ZN(n387) );
  AOI22_X2 U340 ( .A1(\U27/DATA2_29 ), .A2(n871), .B1(\U24/DATA1_29 ), .B2(
        n879), .ZN(n159) );
  AOI22_X2 U341 ( .A1(\U21/DATA1_29 ), .A2(n880), .B1(Diagonal[29]), .B2(n888), 
        .ZN(n160) );
  OAI211_X2 U346 ( .C1(n120), .C2(n911), .A(n157), .B(n158), .ZN(n386) );
  AOI22_X2 U349 ( .A1(\U27/DATA2_30 ), .A2(n871), .B1(\U24/DATA1_30 ), .B2(
        n879), .ZN(n157) );
  AOI22_X2 U351 ( .A1(\U21/DATA1_30 ), .A2(n880), .B1(Diagonal[30]), .B2(n888), 
        .ZN(n158) );
  OAI211_X2 U352 ( .C1(n120), .C2(n910), .A(n155), .B(n156), .ZN(n385) );
  AOI22_X2 U353 ( .A1(\U27/DATA2_31 ), .A2(n871), .B1(\U24/DATA1_31 ), .B2(
        n879), .ZN(n155) );
  AOI22_X2 U354 ( .A1(\U21/DATA1_31 ), .A2(n880), .B1(Diagonal[31]), .B2(n888), 
        .ZN(n156) );
  OAI211_X2 U363 ( .C1(n120), .C2(n909), .A(n153), .B(n154), .ZN(n384) );
  AOI22_X2 U364 ( .A1(\U27/DATA2_32 ), .A2(n871), .B1(\U24/DATA1_32 ), .B2(
        n879), .ZN(n153) );
  AOI22_X2 U365 ( .A1(\U21/DATA1_32 ), .A2(n880), .B1(Diagonal[32]), .B2(n888), 
        .ZN(n154) );
  OAI211_X2 U366 ( .C1(n120), .C2(n908), .A(n151), .B(n152), .ZN(n383) );
  AOI22_X2 U367 ( .A1(\U27/DATA2_33 ), .A2(n871), .B1(\U24/DATA1_33 ), .B2(
        n879), .ZN(n151) );
  AOI22_X2 U368 ( .A1(\U21/DATA1_33 ), .A2(n880), .B1(Diagonal[33]), .B2(n888), 
        .ZN(n152) );
  OAI211_X2 U369 ( .C1(n120), .C2(n907), .A(n149), .B(n150), .ZN(n382) );
  AOI22_X2 U370 ( .A1(\U27/DATA2_34 ), .A2(n871), .B1(\U24/DATA1_34 ), .B2(
        n879), .ZN(n149) );
  AOI22_X2 U371 ( .A1(\U21/DATA1_34 ), .A2(n880), .B1(Diagonal[34]), .B2(n888), 
        .ZN(n150) );
  OAI211_X2 U372 ( .C1(n120), .C2(n906), .A(n147), .B(n148), .ZN(n381) );
  AOI22_X2 U373 ( .A1(\U27/DATA2_35 ), .A2(n871), .B1(\U24/DATA1_35 ), .B2(
        n879), .ZN(n147) );
  AOI22_X2 U374 ( .A1(\U21/DATA1_35 ), .A2(n880), .B1(Diagonal[35]), .B2(n888), 
        .ZN(n148) );
  AOI21_X2 U375 ( .B1(n866), .B2(Element[48]), .A(n347), .ZN(n352) );
  OAI21_X2 U376 ( .B1(\r412/A[0] ), .B2(n891), .A(n882), .ZN(n477) );
  AND2_X4 U377 ( .A1(n247), .A2(n891), .ZN(n223) );
  INV_X4 U378 ( .A(n367), .ZN(n883) );
  INV_X4 U379 ( .A(n368), .ZN(n884) );
  INV_X4 U380 ( .A(n353), .ZN(n885) );
  INV_X4 U381 ( .A(n350), .ZN(n886) );
  INV_X4 U382 ( .A(n348), .ZN(n887) );
  INV_X4 U383 ( .A(n347), .ZN(n888) );
  INV_X4 U384 ( .A(n352), .ZN(n889) );
  INV_X4 U385 ( .A(n364), .ZN(n890) );
  INV_X4 U386 ( .A(n351), .ZN(n891) );
  INV_X4 U387 ( .A(n360), .ZN(n892) );
  INV_X4 U388 ( .A(n357), .ZN(n893) );
  INV_X4 U389 ( .A(\U27/DATA1_47 ), .ZN(n894) );
  INV_X4 U390 ( .A(\U27/DATA1_46 ), .ZN(n895) );
  INV_X4 U391 ( .A(\U27/DATA1_45 ), .ZN(n896) );
  INV_X4 U392 ( .A(\U27/DATA1_44 ), .ZN(n897) );
  INV_X4 U393 ( .A(\U27/DATA1_43 ), .ZN(n898) );
  INV_X4 U394 ( .A(\U27/DATA1_42 ), .ZN(n899) );
  INV_X4 U395 ( .A(\U27/DATA1_41 ), .ZN(n900) );
  INV_X4 U396 ( .A(\U27/DATA1_40 ), .ZN(n901) );
  INV_X4 U397 ( .A(\U27/DATA1_39 ), .ZN(n902) );
  INV_X4 U398 ( .A(\U27/DATA1_38 ), .ZN(n903) );
  INV_X4 U399 ( .A(\U27/DATA1_37 ), .ZN(n904) );
  INV_X4 U400 ( .A(\U27/DATA1_36 ), .ZN(n905) );
  INV_X4 U401 ( .A(\U27/DATA1_35 ), .ZN(n906) );
  INV_X4 U402 ( .A(\U27/DATA1_34 ), .ZN(n907) );
  INV_X4 U403 ( .A(\U27/DATA1_33 ), .ZN(n908) );
  INV_X4 U404 ( .A(\U27/DATA1_32 ), .ZN(n909) );
  INV_X4 U405 ( .A(\U27/DATA1_31 ), .ZN(n910) );
  INV_X4 U406 ( .A(\U27/DATA1_30 ), .ZN(n911) );
  INV_X4 U407 ( .A(\U27/DATA1_29 ), .ZN(n912) );
  INV_X4 U408 ( .A(\U27/DATA1_28 ), .ZN(n913) );
  INV_X4 U409 ( .A(\U27/DATA1_27 ), .ZN(n914) );
  INV_X4 U410 ( .A(\U27/DATA1_26 ), .ZN(n915) );
  INV_X4 U411 ( .A(\U27/DATA1_25 ), .ZN(n916) );
  INV_X4 U412 ( .A(\U27/DATA1_24 ), .ZN(n917) );
  INV_X4 U413 ( .A(\U27/DATA1_23 ), .ZN(n918) );
  INV_X4 U414 ( .A(\U27/DATA1_22 ), .ZN(n919) );
  INV_X4 U415 ( .A(\U27/DATA1_21 ), .ZN(n920) );
  INV_X4 U416 ( .A(\U27/DATA1_20 ), .ZN(n921) );
  INV_X4 U417 ( .A(\U27/DATA1_19 ), .ZN(n922) );
  INV_X4 U418 ( .A(\U27/DATA1_18 ), .ZN(n923) );
  INV_X4 U419 ( .A(\U27/DATA1_17 ), .ZN(n924) );
  INV_X4 U420 ( .A(\U27/DATA1_16 ), .ZN(n925) );
  INV_X4 U421 ( .A(\U27/DATA1_15 ), .ZN(n926) );
  INV_X4 U422 ( .A(\U27/DATA1_14 ), .ZN(n927) );
  INV_X4 U423 ( .A(\U27/DATA1_13 ), .ZN(n928) );
  INV_X4 U424 ( .A(\U27/DATA1_12 ), .ZN(n929) );
  INV_X4 U425 ( .A(\U27/DATA1_11 ), .ZN(n930) );
  INV_X4 U426 ( .A(\U27/DATA1_10 ), .ZN(n931) );
  INV_X4 U427 ( .A(\U27/DATA1_9 ), .ZN(n932) );
  INV_X4 U428 ( .A(\U27/DATA1_8 ), .ZN(n933) );
  INV_X4 U429 ( .A(\U27/DATA1_7 ), .ZN(n934) );
  INV_X4 U430 ( .A(\U27/DATA1_6 ), .ZN(n935) );
  INV_X4 U431 ( .A(\U27/DATA1_5 ), .ZN(n936) );
  INV_X4 U432 ( .A(\U27/DATA1_4 ), .ZN(n937) );
  INV_X4 U433 ( .A(\U27/DATA1_3 ), .ZN(n938) );
  INV_X4 U434 ( .A(\U27/DATA1_2 ), .ZN(n939) );
  INV_X4 U435 ( .A(\U27/DATA1_1 ), .ZN(n940) );
  INV_X4 U436 ( .A(\U27/DATA1_0 ), .ZN(n941) );
  INV_X4 U437 ( .A(\U3/U5/DATA1_2 ), .ZN(n942) );
  INV_X4 U438 ( .A(\U3/U5/DATA1_1 ), .ZN(n943) );
  INV_X4 U439 ( .A(\U3/U5/DATA1_0 ), .ZN(n944) );
  INV_X4 U440 ( .A(\U24/DATA1_47 ), .ZN(n945) );
  INV_X4 U441 ( .A(\U24/DATA1_46 ), .ZN(n946) );
  INV_X4 U442 ( .A(\U24/DATA1_45 ), .ZN(n947) );
  INV_X4 U443 ( .A(\U24/DATA1_44 ), .ZN(n948) );
  INV_X4 U444 ( .A(\U24/DATA1_43 ), .ZN(n949) );
  INV_X4 U445 ( .A(\U24/DATA1_42 ), .ZN(n950) );
  INV_X4 U446 ( .A(\U24/DATA1_41 ), .ZN(n951) );
  INV_X4 U447 ( .A(\U24/DATA1_40 ), .ZN(n952) );
  INV_X4 U448 ( .A(\U24/DATA1_39 ), .ZN(n953) );
  INV_X4 U449 ( .A(\U24/DATA1_38 ), .ZN(n954) );
  INV_X4 U450 ( .A(\U24/DATA1_37 ), .ZN(n955) );
  INV_X4 U451 ( .A(\U24/DATA1_36 ), .ZN(n956) );
  INV_X4 U452 ( .A(\U24/DATA1_35 ), .ZN(n957) );
  INV_X4 U453 ( .A(\U24/DATA1_34 ), .ZN(n958) );
  INV_X4 U454 ( .A(\U24/DATA1_33 ), .ZN(n959) );
  INV_X4 U455 ( .A(\U24/DATA1_32 ), .ZN(n960) );
  INV_X4 U456 ( .A(\U24/DATA1_31 ), .ZN(n961) );
  INV_X4 U457 ( .A(\U24/DATA1_30 ), .ZN(n962) );
  INV_X4 U458 ( .A(\U24/DATA1_29 ), .ZN(n963) );
  INV_X4 U459 ( .A(\U24/DATA1_28 ), .ZN(n964) );
  INV_X4 U460 ( .A(\U24/DATA1_27 ), .ZN(n965) );
  INV_X4 U461 ( .A(\U24/DATA1_26 ), .ZN(n966) );
  INV_X4 U462 ( .A(\U24/DATA1_25 ), .ZN(n967) );
  INV_X4 U463 ( .A(\U24/DATA1_24 ), .ZN(n968) );
  INV_X4 U464 ( .A(\U24/DATA1_23 ), .ZN(n969) );
  INV_X4 U465 ( .A(\U24/DATA1_22 ), .ZN(n970) );
  INV_X4 U466 ( .A(\U24/DATA1_21 ), .ZN(n971) );
  INV_X4 U467 ( .A(\U24/DATA1_20 ), .ZN(n972) );
  INV_X4 U468 ( .A(\U24/DATA1_19 ), .ZN(n973) );
  INV_X4 U469 ( .A(\U24/DATA1_18 ), .ZN(n974) );
  INV_X4 U470 ( .A(\U24/DATA1_17 ), .ZN(n975) );
  INV_X4 U471 ( .A(\U24/DATA1_16 ), .ZN(n976) );
  INV_X4 U472 ( .A(\U24/DATA1_15 ), .ZN(n977) );
  INV_X4 U473 ( .A(\U24/DATA1_14 ), .ZN(n978) );
  INV_X4 U474 ( .A(\U24/DATA1_13 ), .ZN(n979) );
  INV_X4 U475 ( .A(\U24/DATA1_12 ), .ZN(n980) );
  INV_X4 U476 ( .A(\U24/DATA1_11 ), .ZN(n981) );
  INV_X4 U477 ( .A(\U24/DATA1_10 ), .ZN(n982) );
  INV_X4 U478 ( .A(\U24/DATA1_9 ), .ZN(n983) );
  INV_X4 U479 ( .A(\U24/DATA1_8 ), .ZN(n984) );
  INV_X4 U480 ( .A(\U24/DATA1_7 ), .ZN(n985) );
  INV_X4 U481 ( .A(\U24/DATA1_6 ), .ZN(n986) );
  INV_X4 U483 ( .A(\U24/DATA1_5 ), .ZN(n987) );
  INV_X4 U484 ( .A(\U24/DATA1_4 ), .ZN(n988) );
  INV_X4 U485 ( .A(\U24/DATA1_3 ), .ZN(n989) );
  INV_X4 U486 ( .A(\U24/DATA1_2 ), .ZN(n990) );
  INV_X4 U487 ( .A(\U24/DATA1_1 ), .ZN(n991) );
  INV_X4 U488 ( .A(\U24/DATA1_0 ), .ZN(n992) );
  INV_X4 U489 ( .A(\U4/DATA4_3 ), .ZN(n993) );
  INV_X4 U490 ( .A(\U20/DATA1_10 ), .ZN(n994) );
  INV_X4 U491 ( .A(\U20/DATA1_9 ), .ZN(n995) );
  INV_X4 U492 ( .A(\U20/DATA1_8 ), .ZN(n996) );
endmodule


module v_arbiter ( vop1, vop2, vop3, vop4, rowno, clock, Vout, Rowread1, 
        Rowread2, Rowread3, Rowread4, count2 );
  input [47:0] vop1;
  input [47:0] vop2;
  input [47:0] vop3;
  input [47:0] vop4;
  input [10:0] rowno;
  output [47:0] Vout;
  output [8:0] Rowread1;
  output [8:0] Rowread2;
  output [8:0] Rowread3;
  output [8:0] Rowread4;
  input clock, count2;
  wire   \U4/Z_0 , \U4/Z_1 , \U4/Z_2 , \U4/Z_3 , \U4/Z_4 , \U4/Z_5 , \U4/Z_6 ,
         \U4/Z_7 , \U4/Z_8 , \U4/Z_9 , \U4/Z_10 , \U4/Z_11 , \U4/Z_12 ,
         \U4/Z_13 , \U4/Z_14 , \U4/Z_15 , \U4/Z_16 , \U4/Z_17 , \U4/Z_18 ,
         \U4/Z_19 , \U4/Z_20 , \U4/Z_21 , \U4/Z_22 , \U4/Z_23 , \U4/Z_24 ,
         \U4/Z_25 , \U4/Z_26 , \U4/Z_27 , \U4/Z_28 , \U4/Z_29 , \U4/Z_30 ,
         \U4/Z_31 , \U4/Z_32 , \U4/Z_33 , \U4/Z_34 , \U4/Z_35 , \U4/Z_36 ,
         \U4/Z_37 , \U4/Z_38 , \U4/Z_39 , \U4/Z_40 , \U4/Z_41 , \U4/Z_42 ,
         \U4/Z_43 , \U4/Z_44 , \U4/Z_45 , \U4/Z_46 , \U4/Z_47 , \U4/DATA4_0 ,
         \U4/DATA4_1 , \U4/DATA4_2 , \U4/DATA4_3 , \U4/DATA4_4 , \U4/DATA4_5 ,
         \U4/DATA4_6 , \U4/DATA4_7 , \U4/DATA4_8 , \U4/DATA4_9 , \U4/DATA4_10 ,
         \U4/DATA4_11 , \U4/DATA4_12 , \U4/DATA4_13 , \U4/DATA4_14 ,
         \U4/DATA4_15 , \U4/DATA4_16 , \U4/DATA4_17 , \U4/DATA4_18 ,
         \U4/DATA4_19 , \U4/DATA4_20 , \U4/DATA4_21 , \U4/DATA4_22 ,
         \U4/DATA4_23 , \U4/DATA4_24 , \U4/DATA4_25 , \U4/DATA4_26 ,
         \U4/DATA4_27 , \U4/DATA4_28 , \U4/DATA4_29 , \U4/DATA4_30 ,
         \U4/DATA4_31 , \U4/DATA4_32 , \U4/DATA4_33 , \U4/DATA4_34 ,
         \U4/DATA4_35 , \U4/DATA4_36 , \U4/DATA4_37 , \U4/DATA4_38 ,
         \U4/DATA4_39 , \U4/DATA4_40 , \U4/DATA4_41 , \U4/DATA4_42 ,
         \U4/DATA4_43 , \U4/DATA4_44 , \U4/DATA4_45 , \U4/DATA4_46 ,
         \U4/DATA4_47 , \U4/DATA3_0 , \U4/DATA3_1 , \U4/DATA3_2 , \U4/DATA3_3 ,
         \U4/DATA3_4 , \U4/DATA3_5 , \U4/DATA3_6 , \U4/DATA3_7 , \U4/DATA3_8 ,
         \U4/DATA3_9 , \U4/DATA3_10 , \U4/DATA3_11 , \U4/DATA3_12 ,
         \U4/DATA3_13 , \U4/DATA3_14 , \U4/DATA3_15 , \U4/DATA3_16 ,
         \U4/DATA3_17 , \U4/DATA3_18 , \U4/DATA3_19 , \U4/DATA3_20 ,
         \U4/DATA3_21 , \U4/DATA3_22 , \U4/DATA3_23 , \U4/DATA3_24 ,
         \U4/DATA3_25 , \U4/DATA3_26 , \U4/DATA3_27 , \U4/DATA3_28 ,
         \U4/DATA3_29 , \U4/DATA3_30 , \U4/DATA3_31 , \U4/DATA3_32 ,
         \U4/DATA3_33 , \U4/DATA3_34 , \U4/DATA3_35 , \U4/DATA3_36 ,
         \U4/DATA3_37 , \U4/DATA3_38 , \U4/DATA3_39 , \U4/DATA3_40 ,
         \U4/DATA3_41 , \U4/DATA3_42 , \U4/DATA3_43 , \U4/DATA3_44 ,
         \U4/DATA3_45 , \U4/DATA3_46 , \U4/DATA3_47 , \U4/DATA2_0 ,
         \U4/DATA2_1 , \U4/DATA2_2 , \U4/DATA2_3 , \U4/DATA2_4 , \U4/DATA2_5 ,
         \U4/DATA2_6 , \U4/DATA2_7 , \U4/DATA2_8 , \U4/DATA2_9 , \U4/DATA2_10 ,
         \U4/DATA2_11 , \U4/DATA2_12 , \U4/DATA2_13 , \U4/DATA2_14 ,
         \U4/DATA2_15 , \U4/DATA2_16 , \U4/DATA2_17 , \U4/DATA2_18 ,
         \U4/DATA2_19 , \U4/DATA2_20 , \U4/DATA2_21 , \U4/DATA2_22 ,
         \U4/DATA2_23 , \U4/DATA2_24 , \U4/DATA2_25 , \U4/DATA2_26 ,
         \U4/DATA2_27 , \U4/DATA2_28 , \U4/DATA2_29 , \U4/DATA2_30 ,
         \U4/DATA2_31 , \U4/DATA2_32 , \U4/DATA2_33 , \U4/DATA2_34 ,
         \U4/DATA2_35 , \U4/DATA2_36 , \U4/DATA2_37 , \U4/DATA2_38 ,
         \U4/DATA2_39 , \U4/DATA2_40 , \U4/DATA2_41 , \U4/DATA2_42 ,
         \U4/DATA2_43 , \U4/DATA2_44 , \U4/DATA2_45 , \U4/DATA2_46 ,
         \U4/DATA2_47 , \U4/DATA1_0 , \U4/DATA1_1 , \U4/DATA1_2 , \U4/DATA1_3 ,
         \U4/DATA1_4 , \U4/DATA1_5 , \U4/DATA1_6 , \U4/DATA1_7 , \U4/DATA1_8 ,
         \U4/DATA1_9 , \U4/DATA1_10 , \U4/DATA1_11 , \U4/DATA1_12 ,
         \U4/DATA1_13 , \U4/DATA1_14 , \U4/DATA1_15 , \U4/DATA1_16 ,
         \U4/DATA1_17 , \U4/DATA1_18 , \U4/DATA1_19 , \U4/DATA1_20 ,
         \U4/DATA1_21 , \U4/DATA1_22 , \U4/DATA1_23 , \U4/DATA1_24 ,
         \U4/DATA1_25 , \U4/DATA1_26 , \U4/DATA1_27 , \U4/DATA1_28 ,
         \U4/DATA1_29 , \U4/DATA1_30 , \U4/DATA1_31 , \U4/DATA1_32 ,
         \U4/DATA1_33 , \U4/DATA1_34 , \U4/DATA1_35 , \U4/DATA1_36 ,
         \U4/DATA1_37 , \U4/DATA1_38 , \U4/DATA1_39 , \U4/DATA1_40 ,
         \U4/DATA1_41 , \U4/DATA1_42 , \U4/DATA1_43 , \U4/DATA1_44 ,
         \U4/DATA1_45 , \U4/DATA1_46 , \U4/DATA1_47 , \add_29_aco/B[8] ,
         \add_29_aco/A[8] , n2, n3, n5, n6, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n316, n317, n353, n354;
  assign Vout[0] = \U4/Z_0 ;
  assign Vout[1] = \U4/Z_1 ;
  assign Vout[2] = \U4/Z_2 ;
  assign Vout[3] = \U4/Z_3 ;
  assign Vout[4] = \U4/Z_4 ;
  assign Vout[5] = \U4/Z_5 ;
  assign Vout[6] = \U4/Z_6 ;
  assign Vout[7] = \U4/Z_7 ;
  assign Vout[8] = \U4/Z_8 ;
  assign Vout[9] = \U4/Z_9 ;
  assign Vout[10] = \U4/Z_10 ;
  assign Vout[11] = \U4/Z_11 ;
  assign Vout[12] = \U4/Z_12 ;
  assign Vout[13] = \U4/Z_13 ;
  assign Vout[14] = \U4/Z_14 ;
  assign Vout[15] = \U4/Z_15 ;
  assign Vout[16] = \U4/Z_16 ;
  assign Vout[17] = \U4/Z_17 ;
  assign Vout[18] = \U4/Z_18 ;
  assign Vout[19] = \U4/Z_19 ;
  assign Vout[20] = \U4/Z_20 ;
  assign Vout[21] = \U4/Z_21 ;
  assign Vout[22] = \U4/Z_22 ;
  assign Vout[23] = \U4/Z_23 ;
  assign Vout[24] = \U4/Z_24 ;
  assign Vout[25] = \U4/Z_25 ;
  assign Vout[26] = \U4/Z_26 ;
  assign Vout[27] = \U4/Z_27 ;
  assign Vout[28] = \U4/Z_28 ;
  assign Vout[29] = \U4/Z_29 ;
  assign Vout[30] = \U4/Z_30 ;
  assign Vout[31] = \U4/Z_31 ;
  assign Vout[32] = \U4/Z_32 ;
  assign Vout[33] = \U4/Z_33 ;
  assign Vout[34] = \U4/Z_34 ;
  assign Vout[35] = \U4/Z_35 ;
  assign Vout[36] = \U4/Z_36 ;
  assign Vout[37] = \U4/Z_37 ;
  assign Vout[38] = \U4/Z_38 ;
  assign Vout[39] = \U4/Z_39 ;
  assign Vout[40] = \U4/Z_40 ;
  assign Vout[41] = \U4/Z_41 ;
  assign Vout[42] = \U4/Z_42 ;
  assign Vout[43] = \U4/Z_43 ;
  assign Vout[44] = \U4/Z_44 ;
  assign Vout[45] = \U4/Z_45 ;
  assign Vout[46] = \U4/Z_46 ;
  assign Vout[47] = \U4/Z_47 ;
  assign \U4/DATA4_0  = vop4[0];
  assign \U4/DATA4_1  = vop4[1];
  assign \U4/DATA4_2  = vop4[2];
  assign \U4/DATA4_3  = vop4[3];
  assign \U4/DATA4_4  = vop4[4];
  assign \U4/DATA4_5  = vop4[5];
  assign \U4/DATA4_6  = vop4[6];
  assign \U4/DATA4_7  = vop4[7];
  assign \U4/DATA4_8  = vop4[8];
  assign \U4/DATA4_9  = vop4[9];
  assign \U4/DATA4_10  = vop4[10];
  assign \U4/DATA4_11  = vop4[11];
  assign \U4/DATA4_12  = vop4[12];
  assign \U4/DATA4_13  = vop4[13];
  assign \U4/DATA4_14  = vop4[14];
  assign \U4/DATA4_15  = vop4[15];
  assign \U4/DATA4_16  = vop4[16];
  assign \U4/DATA4_17  = vop4[17];
  assign \U4/DATA4_18  = vop4[18];
  assign \U4/DATA4_19  = vop4[19];
  assign \U4/DATA4_20  = vop4[20];
  assign \U4/DATA4_21  = vop4[21];
  assign \U4/DATA4_22  = vop4[22];
  assign \U4/DATA4_23  = vop4[23];
  assign \U4/DATA4_24  = vop4[24];
  assign \U4/DATA4_25  = vop4[25];
  assign \U4/DATA4_26  = vop4[26];
  assign \U4/DATA4_27  = vop4[27];
  assign \U4/DATA4_28  = vop4[28];
  assign \U4/DATA4_29  = vop4[29];
  assign \U4/DATA4_30  = vop4[30];
  assign \U4/DATA4_31  = vop4[31];
  assign \U4/DATA4_32  = vop4[32];
  assign \U4/DATA4_33  = vop4[33];
  assign \U4/DATA4_34  = vop4[34];
  assign \U4/DATA4_35  = vop4[35];
  assign \U4/DATA4_36  = vop4[36];
  assign \U4/DATA4_37  = vop4[37];
  assign \U4/DATA4_38  = vop4[38];
  assign \U4/DATA4_39  = vop4[39];
  assign \U4/DATA4_40  = vop4[40];
  assign \U4/DATA4_41  = vop4[41];
  assign \U4/DATA4_42  = vop4[42];
  assign \U4/DATA4_43  = vop4[43];
  assign \U4/DATA4_44  = vop4[44];
  assign \U4/DATA4_45  = vop4[45];
  assign \U4/DATA4_46  = vop4[46];
  assign \U4/DATA4_47  = vop4[47];
  assign \U4/DATA3_0  = vop3[0];
  assign \U4/DATA3_1  = vop3[1];
  assign \U4/DATA3_2  = vop3[2];
  assign \U4/DATA3_3  = vop3[3];
  assign \U4/DATA3_4  = vop3[4];
  assign \U4/DATA3_5  = vop3[5];
  assign \U4/DATA3_6  = vop3[6];
  assign \U4/DATA3_7  = vop3[7];
  assign \U4/DATA3_8  = vop3[8];
  assign \U4/DATA3_9  = vop3[9];
  assign \U4/DATA3_10  = vop3[10];
  assign \U4/DATA3_11  = vop3[11];
  assign \U4/DATA3_12  = vop3[12];
  assign \U4/DATA3_13  = vop3[13];
  assign \U4/DATA3_14  = vop3[14];
  assign \U4/DATA3_15  = vop3[15];
  assign \U4/DATA3_16  = vop3[16];
  assign \U4/DATA3_17  = vop3[17];
  assign \U4/DATA3_18  = vop3[18];
  assign \U4/DATA3_19  = vop3[19];
  assign \U4/DATA3_20  = vop3[20];
  assign \U4/DATA3_21  = vop3[21];
  assign \U4/DATA3_22  = vop3[22];
  assign \U4/DATA3_23  = vop3[23];
  assign \U4/DATA3_24  = vop3[24];
  assign \U4/DATA3_25  = vop3[25];
  assign \U4/DATA3_26  = vop3[26];
  assign \U4/DATA3_27  = vop3[27];
  assign \U4/DATA3_28  = vop3[28];
  assign \U4/DATA3_29  = vop3[29];
  assign \U4/DATA3_30  = vop3[30];
  assign \U4/DATA3_31  = vop3[31];
  assign \U4/DATA3_32  = vop3[32];
  assign \U4/DATA3_33  = vop3[33];
  assign \U4/DATA3_34  = vop3[34];
  assign \U4/DATA3_35  = vop3[35];
  assign \U4/DATA3_36  = vop3[36];
  assign \U4/DATA3_37  = vop3[37];
  assign \U4/DATA3_38  = vop3[38];
  assign \U4/DATA3_39  = vop3[39];
  assign \U4/DATA3_40  = vop3[40];
  assign \U4/DATA3_41  = vop3[41];
  assign \U4/DATA3_42  = vop3[42];
  assign \U4/DATA3_43  = vop3[43];
  assign \U4/DATA3_44  = vop3[44];
  assign \U4/DATA3_45  = vop3[45];
  assign \U4/DATA3_46  = vop3[46];
  assign \U4/DATA3_47  = vop3[47];
  assign \U4/DATA2_0  = vop2[0];
  assign \U4/DATA2_1  = vop2[1];
  assign \U4/DATA2_2  = vop2[2];
  assign \U4/DATA2_3  = vop2[3];
  assign \U4/DATA2_4  = vop2[4];
  assign \U4/DATA2_5  = vop2[5];
  assign \U4/DATA2_6  = vop2[6];
  assign \U4/DATA2_7  = vop2[7];
  assign \U4/DATA2_8  = vop2[8];
  assign \U4/DATA2_9  = vop2[9];
  assign \U4/DATA2_10  = vop2[10];
  assign \U4/DATA2_11  = vop2[11];
  assign \U4/DATA2_12  = vop2[12];
  assign \U4/DATA2_13  = vop2[13];
  assign \U4/DATA2_14  = vop2[14];
  assign \U4/DATA2_15  = vop2[15];
  assign \U4/DATA2_16  = vop2[16];
  assign \U4/DATA2_17  = vop2[17];
  assign \U4/DATA2_18  = vop2[18];
  assign \U4/DATA2_19  = vop2[19];
  assign \U4/DATA2_20  = vop2[20];
  assign \U4/DATA2_21  = vop2[21];
  assign \U4/DATA2_22  = vop2[22];
  assign \U4/DATA2_23  = vop2[23];
  assign \U4/DATA2_24  = vop2[24];
  assign \U4/DATA2_25  = vop2[25];
  assign \U4/DATA2_26  = vop2[26];
  assign \U4/DATA2_27  = vop2[27];
  assign \U4/DATA2_28  = vop2[28];
  assign \U4/DATA2_29  = vop2[29];
  assign \U4/DATA2_30  = vop2[30];
  assign \U4/DATA2_31  = vop2[31];
  assign \U4/DATA2_32  = vop2[32];
  assign \U4/DATA2_33  = vop2[33];
  assign \U4/DATA2_34  = vop2[34];
  assign \U4/DATA2_35  = vop2[35];
  assign \U4/DATA2_36  = vop2[36];
  assign \U4/DATA2_37  = vop2[37];
  assign \U4/DATA2_38  = vop2[38];
  assign \U4/DATA2_39  = vop2[39];
  assign \U4/DATA2_40  = vop2[40];
  assign \U4/DATA2_41  = vop2[41];
  assign \U4/DATA2_42  = vop2[42];
  assign \U4/DATA2_43  = vop2[43];
  assign \U4/DATA2_44  = vop2[44];
  assign \U4/DATA2_45  = vop2[45];
  assign \U4/DATA2_46  = vop2[46];
  assign \U4/DATA2_47  = vop2[47];
  assign \U4/DATA1_0  = vop1[0];
  assign \U4/DATA1_1  = vop1[1];
  assign \U4/DATA1_2  = vop1[2];
  assign \U4/DATA1_3  = vop1[3];
  assign \U4/DATA1_4  = vop1[4];
  assign \U4/DATA1_5  = vop1[5];
  assign \U4/DATA1_6  = vop1[6];
  assign \U4/DATA1_7  = vop1[7];
  assign \U4/DATA1_8  = vop1[8];
  assign \U4/DATA1_9  = vop1[9];
  assign \U4/DATA1_10  = vop1[10];
  assign \U4/DATA1_11  = vop1[11];
  assign \U4/DATA1_12  = vop1[12];
  assign \U4/DATA1_13  = vop1[13];
  assign \U4/DATA1_14  = vop1[14];
  assign \U4/DATA1_15  = vop1[15];
  assign \U4/DATA1_16  = vop1[16];
  assign \U4/DATA1_17  = vop1[17];
  assign \U4/DATA1_18  = vop1[18];
  assign \U4/DATA1_19  = vop1[19];
  assign \U4/DATA1_20  = vop1[20];
  assign \U4/DATA1_21  = vop1[21];
  assign \U4/DATA1_22  = vop1[22];
  assign \U4/DATA1_23  = vop1[23];
  assign \U4/DATA1_24  = vop1[24];
  assign \U4/DATA1_25  = vop1[25];
  assign \U4/DATA1_26  = vop1[26];
  assign \U4/DATA1_27  = vop1[27];
  assign \U4/DATA1_28  = vop1[28];
  assign \U4/DATA1_29  = vop1[29];
  assign \U4/DATA1_30  = vop1[30];
  assign \U4/DATA1_31  = vop1[31];
  assign \U4/DATA1_32  = vop1[32];
  assign \U4/DATA1_33  = vop1[33];
  assign \U4/DATA1_34  = vop1[34];
  assign \U4/DATA1_35  = vop1[35];
  assign \U4/DATA1_36  = vop1[36];
  assign \U4/DATA1_37  = vop1[37];
  assign \U4/DATA1_38  = vop1[38];
  assign \U4/DATA1_39  = vop1[39];
  assign \U4/DATA1_40  = vop1[40];
  assign \U4/DATA1_41  = vop1[41];
  assign \U4/DATA1_42  = vop1[42];
  assign \U4/DATA1_43  = vop1[43];
  assign \U4/DATA1_44  = vop1[44];
  assign \U4/DATA1_45  = vop1[45];
  assign \U4/DATA1_46  = vop1[46];
  assign \U4/DATA1_47  = vop1[47];
  assign \add_29_aco/B[8]  = count2;
  assign \add_29_aco/A[8]  = rowno[10];

  NAND2_X2 U2 ( .A1(n2), .A2(n3), .ZN(\U4/Z_9 ) );
  NAND2_X2 U5 ( .A1(n8), .A2(n9), .ZN(\U4/Z_8 ) );
  NAND2_X2 U8 ( .A1(n10), .A2(n11), .ZN(\U4/Z_7 ) );
  NAND2_X2 U11 ( .A1(n12), .A2(n13), .ZN(\U4/Z_6 ) );
  NAND2_X2 U14 ( .A1(n14), .A2(n15), .ZN(\U4/Z_5 ) );
  NAND2_X2 U17 ( .A1(n16), .A2(n17), .ZN(\U4/Z_47 ) );
  NAND2_X2 U20 ( .A1(n18), .A2(n19), .ZN(\U4/Z_46 ) );
  NAND2_X2 U23 ( .A1(n20), .A2(n21), .ZN(\U4/Z_45 ) );
  NAND2_X2 U26 ( .A1(n22), .A2(n23), .ZN(\U4/Z_44 ) );
  NAND2_X2 U29 ( .A1(n24), .A2(n25), .ZN(\U4/Z_43 ) );
  NAND2_X2 U32 ( .A1(n26), .A2(n27), .ZN(\U4/Z_42 ) );
  NAND2_X2 U35 ( .A1(n28), .A2(n29), .ZN(\U4/Z_41 ) );
  NAND2_X2 U38 ( .A1(n30), .A2(n31), .ZN(\U4/Z_40 ) );
  NAND2_X2 U41 ( .A1(n32), .A2(n33), .ZN(\U4/Z_4 ) );
  NAND2_X2 U44 ( .A1(n34), .A2(n35), .ZN(\U4/Z_39 ) );
  NAND2_X2 U47 ( .A1(n36), .A2(n37), .ZN(\U4/Z_38 ) );
  NAND2_X2 U50 ( .A1(n38), .A2(n39), .ZN(\U4/Z_37 ) );
  NAND2_X2 U53 ( .A1(n40), .A2(n41), .ZN(\U4/Z_36 ) );
  NAND2_X2 U56 ( .A1(n42), .A2(n43), .ZN(\U4/Z_35 ) );
  NAND2_X2 U59 ( .A1(n44), .A2(n45), .ZN(\U4/Z_34 ) );
  NAND2_X2 U62 ( .A1(n46), .A2(n47), .ZN(\U4/Z_33 ) );
  NAND2_X2 U65 ( .A1(n48), .A2(n49), .ZN(\U4/Z_32 ) );
  NAND2_X2 U68 ( .A1(n50), .A2(n51), .ZN(\U4/Z_31 ) );
  NAND2_X2 U71 ( .A1(n52), .A2(n53), .ZN(\U4/Z_30 ) );
  NAND2_X2 U74 ( .A1(n54), .A2(n55), .ZN(\U4/Z_3 ) );
  NAND2_X2 U77 ( .A1(n56), .A2(n57), .ZN(\U4/Z_29 ) );
  NAND2_X2 U80 ( .A1(n58), .A2(n59), .ZN(\U4/Z_28 ) );
  NAND2_X2 U83 ( .A1(n60), .A2(n61), .ZN(\U4/Z_27 ) );
  NAND2_X2 U86 ( .A1(n62), .A2(n63), .ZN(\U4/Z_26 ) );
  NAND2_X2 U89 ( .A1(n64), .A2(n65), .ZN(\U4/Z_25 ) );
  NAND2_X2 U92 ( .A1(n66), .A2(n67), .ZN(\U4/Z_24 ) );
  NAND2_X2 U95 ( .A1(n68), .A2(n69), .ZN(\U4/Z_23 ) );
  NAND2_X2 U98 ( .A1(n70), .A2(n71), .ZN(\U4/Z_22 ) );
  NAND2_X2 U101 ( .A1(n72), .A2(n73), .ZN(\U4/Z_21 ) );
  NAND2_X2 U104 ( .A1(n74), .A2(n75), .ZN(\U4/Z_20 ) );
  NAND2_X2 U107 ( .A1(n76), .A2(n77), .ZN(\U4/Z_2 ) );
  NAND2_X2 U110 ( .A1(n78), .A2(n79), .ZN(\U4/Z_19 ) );
  NAND2_X2 U113 ( .A1(n80), .A2(n81), .ZN(\U4/Z_18 ) );
  NAND2_X2 U116 ( .A1(n82), .A2(n83), .ZN(\U4/Z_17 ) );
  NAND2_X2 U119 ( .A1(n84), .A2(n85), .ZN(\U4/Z_16 ) );
  NAND2_X2 U122 ( .A1(n86), .A2(n87), .ZN(\U4/Z_15 ) );
  NAND2_X2 U125 ( .A1(n88), .A2(n89), .ZN(\U4/Z_14 ) );
  NAND2_X2 U128 ( .A1(n90), .A2(n91), .ZN(\U4/Z_13 ) );
  NAND2_X2 U131 ( .A1(n92), .A2(n93), .ZN(\U4/Z_12 ) );
  NAND2_X2 U134 ( .A1(n94), .A2(n95), .ZN(\U4/Z_11 ) );
  NAND2_X2 U137 ( .A1(n96), .A2(n97), .ZN(\U4/Z_10 ) );
  NAND2_X2 U140 ( .A1(n98), .A2(n99), .ZN(\U4/Z_1 ) );
  NAND2_X2 U143 ( .A1(n100), .A2(n101), .ZN(\U4/Z_0 ) );
  NOR2_X4 U3 ( .A1(rowno[1]), .A2(rowno[0]), .ZN(n316) );
  NOR2_X4 U4 ( .A1(n354), .A2(rowno[1]), .ZN(n6) );
  AND2_X4 U6 ( .A1(rowno[1]), .A2(rowno[0]), .ZN(n317) );
  AND2_X4 U7 ( .A1(rowno[1]), .A2(n354), .ZN(n5) );
  BUF_X4 U9 ( .A(Rowread3[8]), .Z(Rowread4[8]) );
  BUF_X4 U10 ( .A(Rowread3[8]), .Z(Rowread2[8]) );
  BUF_X4 U12 ( .A(Rowread3[8]), .Z(Rowread1[8]) );
  AOI22_X2 U13 ( .A1(\U4/DATA2_0 ), .A2(n6), .B1(\U4/DATA1_0 ), .B2(n316), 
        .ZN(n100) );
  AOI22_X2 U15 ( .A1(\U4/DATA4_0 ), .A2(n317), .B1(\U4/DATA3_0 ), .B2(n5), 
        .ZN(n101) );
  AOI22_X2 U16 ( .A1(\U4/DATA2_1 ), .A2(n6), .B1(\U4/DATA1_1 ), .B2(n316), 
        .ZN(n98) );
  AOI22_X2 U18 ( .A1(\U4/DATA4_1 ), .A2(n317), .B1(\U4/DATA3_1 ), .B2(n5), 
        .ZN(n99) );
  AOI22_X2 U19 ( .A1(\U4/DATA2_2 ), .A2(n6), .B1(\U4/DATA1_2 ), .B2(n316), 
        .ZN(n76) );
  AOI22_X2 U21 ( .A1(\U4/DATA4_2 ), .A2(n317), .B1(\U4/DATA3_2 ), .B2(n5), 
        .ZN(n77) );
  AOI22_X2 U22 ( .A1(\U4/DATA2_3 ), .A2(n6), .B1(\U4/DATA1_3 ), .B2(n316), 
        .ZN(n54) );
  AOI22_X2 U24 ( .A1(\U4/DATA4_3 ), .A2(n317), .B1(\U4/DATA3_3 ), .B2(n5), 
        .ZN(n55) );
  AOI22_X2 U25 ( .A1(\U4/DATA2_4 ), .A2(n6), .B1(\U4/DATA1_4 ), .B2(n316), 
        .ZN(n32) );
  AOI22_X2 U27 ( .A1(\U4/DATA4_4 ), .A2(n317), .B1(\U4/DATA3_4 ), .B2(n5), 
        .ZN(n33) );
  AOI22_X2 U28 ( .A1(\U4/DATA2_5 ), .A2(n6), .B1(\U4/DATA1_5 ), .B2(n316), 
        .ZN(n14) );
  AOI22_X2 U30 ( .A1(\U4/DATA4_5 ), .A2(n317), .B1(\U4/DATA3_5 ), .B2(n5), 
        .ZN(n15) );
  AOI22_X2 U31 ( .A1(\U4/DATA2_6 ), .A2(n6), .B1(\U4/DATA1_6 ), .B2(n316), 
        .ZN(n12) );
  AOI22_X2 U33 ( .A1(\U4/DATA4_6 ), .A2(n317), .B1(\U4/DATA3_6 ), .B2(n5), 
        .ZN(n13) );
  AOI22_X2 U34 ( .A1(\U4/DATA2_7 ), .A2(n6), .B1(\U4/DATA1_7 ), .B2(n316), 
        .ZN(n10) );
  AOI22_X2 U36 ( .A1(\U4/DATA4_7 ), .A2(n317), .B1(\U4/DATA3_7 ), .B2(n5), 
        .ZN(n11) );
  AOI22_X2 U37 ( .A1(\U4/DATA2_8 ), .A2(n6), .B1(\U4/DATA1_8 ), .B2(n316), 
        .ZN(n8) );
  AOI22_X2 U39 ( .A1(\U4/DATA4_8 ), .A2(n317), .B1(\U4/DATA3_8 ), .B2(n5), 
        .ZN(n9) );
  AOI22_X2 U40 ( .A1(\U4/DATA2_9 ), .A2(n6), .B1(\U4/DATA1_9 ), .B2(n316), 
        .ZN(n2) );
  AOI22_X2 U42 ( .A1(\U4/DATA4_9 ), .A2(n317), .B1(\U4/DATA3_9 ), .B2(n5), 
        .ZN(n3) );
  AOI22_X2 U43 ( .A1(\U4/DATA2_10 ), .A2(n6), .B1(\U4/DATA1_10 ), .B2(n316), 
        .ZN(n96) );
  AOI22_X2 U45 ( .A1(\U4/DATA4_10 ), .A2(n317), .B1(\U4/DATA3_10 ), .B2(n5), 
        .ZN(n97) );
  AOI22_X2 U46 ( .A1(\U4/DATA2_11 ), .A2(n6), .B1(\U4/DATA1_11 ), .B2(n316), 
        .ZN(n94) );
  AOI22_X2 U48 ( .A1(\U4/DATA4_11 ), .A2(n317), .B1(\U4/DATA3_11 ), .B2(n5), 
        .ZN(n95) );
  AOI22_X2 U49 ( .A1(\U4/DATA2_12 ), .A2(n6), .B1(\U4/DATA1_12 ), .B2(n316), 
        .ZN(n92) );
  AOI22_X2 U51 ( .A1(\U4/DATA4_12 ), .A2(n317), .B1(\U4/DATA3_12 ), .B2(n5), 
        .ZN(n93) );
  AOI22_X2 U52 ( .A1(\U4/DATA2_13 ), .A2(n6), .B1(\U4/DATA1_13 ), .B2(n316), 
        .ZN(n90) );
  AOI22_X2 U54 ( .A1(\U4/DATA4_13 ), .A2(n317), .B1(\U4/DATA3_13 ), .B2(n5), 
        .ZN(n91) );
  AOI22_X2 U55 ( .A1(\U4/DATA2_14 ), .A2(n6), .B1(\U4/DATA1_14 ), .B2(n316), 
        .ZN(n88) );
  AOI22_X2 U57 ( .A1(\U4/DATA4_14 ), .A2(n317), .B1(\U4/DATA3_14 ), .B2(n5), 
        .ZN(n89) );
  AOI22_X2 U58 ( .A1(\U4/DATA2_15 ), .A2(n6), .B1(\U4/DATA1_15 ), .B2(n316), 
        .ZN(n86) );
  AOI22_X2 U60 ( .A1(\U4/DATA4_15 ), .A2(n317), .B1(\U4/DATA3_15 ), .B2(n5), 
        .ZN(n87) );
  AOI22_X2 U61 ( .A1(\U4/DATA2_16 ), .A2(n6), .B1(\U4/DATA1_16 ), .B2(n316), 
        .ZN(n84) );
  AOI22_X2 U63 ( .A1(\U4/DATA4_16 ), .A2(n317), .B1(\U4/DATA3_16 ), .B2(n5), 
        .ZN(n85) );
  AOI22_X2 U64 ( .A1(\U4/DATA2_17 ), .A2(n6), .B1(\U4/DATA1_17 ), .B2(n316), 
        .ZN(n82) );
  AOI22_X2 U66 ( .A1(\U4/DATA4_17 ), .A2(n317), .B1(\U4/DATA3_17 ), .B2(n5), 
        .ZN(n83) );
  AOI22_X2 U67 ( .A1(\U4/DATA2_18 ), .A2(n6), .B1(\U4/DATA1_18 ), .B2(n316), 
        .ZN(n80) );
  AOI22_X2 U69 ( .A1(\U4/DATA4_18 ), .A2(n317), .B1(\U4/DATA3_18 ), .B2(n5), 
        .ZN(n81) );
  AOI22_X2 U70 ( .A1(\U4/DATA2_19 ), .A2(n6), .B1(\U4/DATA1_19 ), .B2(n316), 
        .ZN(n78) );
  AOI22_X2 U72 ( .A1(\U4/DATA4_19 ), .A2(n317), .B1(\U4/DATA3_19 ), .B2(n5), 
        .ZN(n79) );
  AOI22_X2 U73 ( .A1(\U4/DATA2_20 ), .A2(n6), .B1(\U4/DATA1_20 ), .B2(n316), 
        .ZN(n74) );
  AOI22_X2 U75 ( .A1(\U4/DATA4_20 ), .A2(n317), .B1(\U4/DATA3_20 ), .B2(n5), 
        .ZN(n75) );
  AOI22_X2 U76 ( .A1(\U4/DATA2_21 ), .A2(n6), .B1(\U4/DATA1_21 ), .B2(n316), 
        .ZN(n72) );
  AOI22_X2 U78 ( .A1(\U4/DATA4_21 ), .A2(n317), .B1(\U4/DATA3_21 ), .B2(n5), 
        .ZN(n73) );
  AOI22_X2 U79 ( .A1(\U4/DATA2_22 ), .A2(n6), .B1(\U4/DATA1_22 ), .B2(n316), 
        .ZN(n70) );
  AOI22_X2 U81 ( .A1(\U4/DATA4_22 ), .A2(n317), .B1(\U4/DATA3_22 ), .B2(n5), 
        .ZN(n71) );
  AOI22_X2 U82 ( .A1(\U4/DATA2_23 ), .A2(n6), .B1(\U4/DATA1_23 ), .B2(n316), 
        .ZN(n68) );
  AOI22_X2 U84 ( .A1(\U4/DATA4_23 ), .A2(n317), .B1(\U4/DATA3_23 ), .B2(n5), 
        .ZN(n69) );
  AOI22_X2 U85 ( .A1(\U4/DATA2_24 ), .A2(n6), .B1(\U4/DATA1_24 ), .B2(n316), 
        .ZN(n66) );
  AOI22_X2 U87 ( .A1(\U4/DATA4_24 ), .A2(n317), .B1(\U4/DATA3_24 ), .B2(n5), 
        .ZN(n67) );
  AOI22_X2 U88 ( .A1(\U4/DATA2_25 ), .A2(n6), .B1(\U4/DATA1_25 ), .B2(n316), 
        .ZN(n64) );
  AOI22_X2 U90 ( .A1(\U4/DATA4_25 ), .A2(n317), .B1(\U4/DATA3_25 ), .B2(n5), 
        .ZN(n65) );
  AOI22_X2 U91 ( .A1(\U4/DATA2_26 ), .A2(n6), .B1(\U4/DATA1_26 ), .B2(n316), 
        .ZN(n62) );
  AOI22_X2 U93 ( .A1(\U4/DATA4_26 ), .A2(n317), .B1(\U4/DATA3_26 ), .B2(n5), 
        .ZN(n63) );
  AOI22_X2 U94 ( .A1(\U4/DATA2_27 ), .A2(n6), .B1(\U4/DATA1_27 ), .B2(n316), 
        .ZN(n60) );
  AOI22_X2 U96 ( .A1(\U4/DATA4_27 ), .A2(n317), .B1(\U4/DATA3_27 ), .B2(n5), 
        .ZN(n61) );
  AOI22_X2 U97 ( .A1(\U4/DATA2_28 ), .A2(n6), .B1(\U4/DATA1_28 ), .B2(n316), 
        .ZN(n58) );
  AOI22_X2 U99 ( .A1(\U4/DATA4_28 ), .A2(n317), .B1(\U4/DATA3_28 ), .B2(n5), 
        .ZN(n59) );
  AOI22_X2 U100 ( .A1(\U4/DATA2_29 ), .A2(n6), .B1(\U4/DATA1_29 ), .B2(n316), 
        .ZN(n56) );
  AOI22_X2 U102 ( .A1(\U4/DATA4_29 ), .A2(n317), .B1(\U4/DATA3_29 ), .B2(n5), 
        .ZN(n57) );
  AOI22_X2 U103 ( .A1(\U4/DATA2_30 ), .A2(n6), .B1(\U4/DATA1_30 ), .B2(n316), 
        .ZN(n52) );
  AOI22_X2 U105 ( .A1(\U4/DATA4_30 ), .A2(n317), .B1(\U4/DATA3_30 ), .B2(n5), 
        .ZN(n53) );
  AOI22_X2 U106 ( .A1(\U4/DATA2_31 ), .A2(n6), .B1(\U4/DATA1_31 ), .B2(n316), 
        .ZN(n50) );
  AOI22_X2 U108 ( .A1(\U4/DATA4_31 ), .A2(n317), .B1(\U4/DATA3_31 ), .B2(n5), 
        .ZN(n51) );
  AOI22_X2 U109 ( .A1(\U4/DATA2_32 ), .A2(n6), .B1(\U4/DATA1_32 ), .B2(n316), 
        .ZN(n48) );
  AOI22_X2 U111 ( .A1(\U4/DATA4_32 ), .A2(n317), .B1(\U4/DATA3_32 ), .B2(n5), 
        .ZN(n49) );
  AOI22_X2 U112 ( .A1(\U4/DATA2_33 ), .A2(n6), .B1(\U4/DATA1_33 ), .B2(n316), 
        .ZN(n46) );
  AOI22_X2 U114 ( .A1(\U4/DATA4_33 ), .A2(n317), .B1(\U4/DATA3_33 ), .B2(n5), 
        .ZN(n47) );
  AOI22_X2 U115 ( .A1(\U4/DATA2_34 ), .A2(n6), .B1(\U4/DATA1_34 ), .B2(n316), 
        .ZN(n44) );
  AOI22_X2 U117 ( .A1(\U4/DATA4_34 ), .A2(n317), .B1(\U4/DATA3_34 ), .B2(n5), 
        .ZN(n45) );
  AOI22_X2 U118 ( .A1(\U4/DATA2_35 ), .A2(n6), .B1(\U4/DATA1_35 ), .B2(n316), 
        .ZN(n42) );
  AOI22_X2 U120 ( .A1(\U4/DATA4_35 ), .A2(n317), .B1(\U4/DATA3_35 ), .B2(n5), 
        .ZN(n43) );
  AOI22_X2 U121 ( .A1(\U4/DATA2_36 ), .A2(n6), .B1(\U4/DATA1_36 ), .B2(n316), 
        .ZN(n40) );
  AOI22_X2 U123 ( .A1(\U4/DATA4_36 ), .A2(n317), .B1(\U4/DATA3_36 ), .B2(n5), 
        .ZN(n41) );
  AOI22_X2 U124 ( .A1(\U4/DATA2_37 ), .A2(n6), .B1(\U4/DATA1_37 ), .B2(n316), 
        .ZN(n38) );
  AOI22_X2 U126 ( .A1(\U4/DATA4_37 ), .A2(n317), .B1(\U4/DATA3_37 ), .B2(n5), 
        .ZN(n39) );
  AOI22_X2 U127 ( .A1(\U4/DATA2_38 ), .A2(n6), .B1(\U4/DATA1_38 ), .B2(n316), 
        .ZN(n36) );
  AOI22_X2 U129 ( .A1(\U4/DATA4_38 ), .A2(n317), .B1(\U4/DATA3_38 ), .B2(n5), 
        .ZN(n37) );
  AOI22_X2 U130 ( .A1(\U4/DATA2_39 ), .A2(n6), .B1(\U4/DATA1_39 ), .B2(n316), 
        .ZN(n34) );
  AOI22_X2 U132 ( .A1(\U4/DATA4_39 ), .A2(n317), .B1(\U4/DATA3_39 ), .B2(n5), 
        .ZN(n35) );
  AOI22_X2 U133 ( .A1(\U4/DATA2_40 ), .A2(n6), .B1(\U4/DATA1_40 ), .B2(n316), 
        .ZN(n30) );
  AOI22_X2 U135 ( .A1(\U4/DATA4_40 ), .A2(n317), .B1(\U4/DATA3_40 ), .B2(n5), 
        .ZN(n31) );
  AOI22_X2 U136 ( .A1(\U4/DATA2_41 ), .A2(n6), .B1(\U4/DATA1_41 ), .B2(n316), 
        .ZN(n28) );
  AOI22_X2 U138 ( .A1(\U4/DATA4_41 ), .A2(n317), .B1(\U4/DATA3_41 ), .B2(n5), 
        .ZN(n29) );
  AOI22_X2 U139 ( .A1(\U4/DATA2_42 ), .A2(n6), .B1(\U4/DATA1_42 ), .B2(n316), 
        .ZN(n26) );
  AOI22_X2 U141 ( .A1(\U4/DATA4_42 ), .A2(n317), .B1(\U4/DATA3_42 ), .B2(n5), 
        .ZN(n27) );
  AOI22_X2 U142 ( .A1(\U4/DATA2_43 ), .A2(n6), .B1(\U4/DATA1_43 ), .B2(n316), 
        .ZN(n24) );
  AOI22_X2 U144 ( .A1(\U4/DATA4_43 ), .A2(n317), .B1(\U4/DATA3_43 ), .B2(n5), 
        .ZN(n25) );
  AOI22_X2 U145 ( .A1(\U4/DATA2_44 ), .A2(n6), .B1(\U4/DATA1_44 ), .B2(n316), 
        .ZN(n22) );
  AOI22_X2 U146 ( .A1(\U4/DATA4_44 ), .A2(n317), .B1(\U4/DATA3_44 ), .B2(n5), 
        .ZN(n23) );
  AOI22_X2 U147 ( .A1(\U4/DATA2_45 ), .A2(n6), .B1(\U4/DATA1_45 ), .B2(n316), 
        .ZN(n20) );
  AOI22_X2 U148 ( .A1(\U4/DATA4_45 ), .A2(n317), .B1(\U4/DATA3_45 ), .B2(n5), 
        .ZN(n21) );
  AOI22_X2 U149 ( .A1(\U4/DATA2_46 ), .A2(n6), .B1(\U4/DATA1_46 ), .B2(n316), 
        .ZN(n18) );
  AOI22_X2 U150 ( .A1(\U4/DATA4_46 ), .A2(n317), .B1(\U4/DATA3_46 ), .B2(n5), 
        .ZN(n19) );
  AOI22_X2 U151 ( .A1(\U4/DATA2_47 ), .A2(n6), .B1(\U4/DATA1_47 ), .B2(n316), 
        .ZN(n16) );
  AOI22_X2 U152 ( .A1(\U4/DATA4_47 ), .A2(n317), .B1(\U4/DATA3_47 ), .B2(n5), 
        .ZN(n17) );
  BUF_X4 U153 ( .A(rowno[3]), .Z(Rowread4[1]) );
  BUF_X4 U154 ( .A(rowno[4]), .Z(Rowread4[2]) );
  BUF_X4 U155 ( .A(rowno[5]), .Z(Rowread4[3]) );
  BUF_X4 U156 ( .A(rowno[6]), .Z(Rowread4[4]) );
  BUF_X4 U157 ( .A(rowno[7]), .Z(Rowread4[5]) );
  BUF_X4 U158 ( .A(rowno[8]), .Z(Rowread4[6]) );
  BUF_X4 U159 ( .A(rowno[9]), .Z(Rowread4[7]) );
  BUF_X4 U160 ( .A(rowno[3]), .Z(Rowread3[1]) );
  BUF_X4 U161 ( .A(rowno[4]), .Z(Rowread3[2]) );
  BUF_X4 U162 ( .A(rowno[5]), .Z(Rowread3[3]) );
  BUF_X4 U163 ( .A(rowno[6]), .Z(Rowread3[4]) );
  BUF_X4 U164 ( .A(rowno[7]), .Z(Rowread3[5]) );
  BUF_X4 U165 ( .A(rowno[8]), .Z(Rowread3[6]) );
  BUF_X4 U166 ( .A(rowno[9]), .Z(Rowread3[7]) );
  BUF_X4 U167 ( .A(rowno[3]), .Z(Rowread2[1]) );
  BUF_X4 U168 ( .A(rowno[4]), .Z(Rowread2[2]) );
  BUF_X4 U169 ( .A(rowno[5]), .Z(Rowread2[3]) );
  BUF_X4 U170 ( .A(rowno[6]), .Z(Rowread2[4]) );
  BUF_X4 U171 ( .A(rowno[7]), .Z(Rowread2[5]) );
  BUF_X4 U172 ( .A(rowno[8]), .Z(Rowread2[6]) );
  BUF_X4 U173 ( .A(rowno[9]), .Z(Rowread2[7]) );
  BUF_X4 U174 ( .A(rowno[3]), .Z(Rowread1[1]) );
  BUF_X4 U175 ( .A(rowno[4]), .Z(Rowread1[2]) );
  BUF_X4 U176 ( .A(rowno[5]), .Z(Rowread1[3]) );
  BUF_X4 U177 ( .A(rowno[6]), .Z(Rowread1[4]) );
  BUF_X4 U178 ( .A(rowno[7]), .Z(Rowread1[5]) );
  BUF_X4 U179 ( .A(rowno[8]), .Z(Rowread1[6]) );
  BUF_X4 U180 ( .A(rowno[9]), .Z(Rowread1[7]) );
  BUF_X4 U181 ( .A(rowno[2]), .Z(Rowread3[0]) );
  BUF_X4 U182 ( .A(rowno[2]), .Z(Rowread2[0]) );
  BUF_X4 U183 ( .A(rowno[2]), .Z(Rowread1[0]) );
  BUF_X4 U184 ( .A(rowno[2]), .Z(Rowread4[0]) );
  XNOR2_X2 U185 ( .A(\add_29_aco/B[8] ), .B(n353), .ZN(Rowread3[8]) );
  INV_X4 U186 ( .A(\add_29_aco/A[8] ), .ZN(n353) );
  INV_X4 U187 ( .A(rowno[0]), .ZN(n354) );
endmodule


module sync ( clock, ElementY, ElementV, SyncY, SyncV );
  input [48:0] ElementY;
  input [47:0] ElementV;
  output [48:0] SyncY;
  output [47:0] SyncV;
  input clock;


  DFF_X1 \SyncY_reg[48]  ( .D(ElementY[48]), .CK(clock), .Q(SyncY[48]) );
  DFF_X1 \SyncY_reg[47]  ( .D(ElementY[47]), .CK(clock), .Q(SyncY[47]) );
  DFF_X1 \SyncY_reg[46]  ( .D(ElementY[46]), .CK(clock), .Q(SyncY[46]) );
  DFF_X1 \SyncY_reg[45]  ( .D(ElementY[45]), .CK(clock), .Q(SyncY[45]) );
  DFF_X1 \SyncY_reg[44]  ( .D(ElementY[44]), .CK(clock), .Q(SyncY[44]) );
  DFF_X1 \SyncY_reg[43]  ( .D(ElementY[43]), .CK(clock), .Q(SyncY[43]) );
  DFF_X1 \SyncY_reg[42]  ( .D(ElementY[42]), .CK(clock), .Q(SyncY[42]) );
  DFF_X1 \SyncY_reg[41]  ( .D(ElementY[41]), .CK(clock), .Q(SyncY[41]) );
  DFF_X1 \SyncY_reg[40]  ( .D(ElementY[40]), .CK(clock), .Q(SyncY[40]) );
  DFF_X1 \SyncY_reg[39]  ( .D(ElementY[39]), .CK(clock), .Q(SyncY[39]) );
  DFF_X1 \SyncY_reg[38]  ( .D(ElementY[38]), .CK(clock), .Q(SyncY[38]) );
  DFF_X1 \SyncY_reg[37]  ( .D(ElementY[37]), .CK(clock), .Q(SyncY[37]) );
  DFF_X1 \SyncY_reg[36]  ( .D(ElementY[36]), .CK(clock), .Q(SyncY[36]) );
  DFF_X1 \SyncY_reg[35]  ( .D(ElementY[35]), .CK(clock), .Q(SyncY[35]) );
  DFF_X1 \SyncY_reg[34]  ( .D(ElementY[34]), .CK(clock), .Q(SyncY[34]) );
  DFF_X1 \SyncY_reg[33]  ( .D(ElementY[33]), .CK(clock), .Q(SyncY[33]) );
  DFF_X1 \SyncY_reg[32]  ( .D(ElementY[32]), .CK(clock), .Q(SyncY[32]) );
  DFF_X1 \SyncY_reg[31]  ( .D(ElementY[31]), .CK(clock), .Q(SyncY[31]) );
  DFF_X1 \SyncY_reg[30]  ( .D(ElementY[30]), .CK(clock), .Q(SyncY[30]) );
  DFF_X1 \SyncY_reg[29]  ( .D(ElementY[29]), .CK(clock), .Q(SyncY[29]) );
  DFF_X1 \SyncY_reg[28]  ( .D(ElementY[28]), .CK(clock), .Q(SyncY[28]) );
  DFF_X1 \SyncY_reg[27]  ( .D(ElementY[27]), .CK(clock), .Q(SyncY[27]) );
  DFF_X1 \SyncY_reg[26]  ( .D(ElementY[26]), .CK(clock), .Q(SyncY[26]) );
  DFF_X1 \SyncY_reg[25]  ( .D(ElementY[25]), .CK(clock), .Q(SyncY[25]) );
  DFF_X1 \SyncY_reg[24]  ( .D(ElementY[24]), .CK(clock), .Q(SyncY[24]) );
  DFF_X1 \SyncY_reg[23]  ( .D(ElementY[23]), .CK(clock), .Q(SyncY[23]) );
  DFF_X1 \SyncY_reg[22]  ( .D(ElementY[22]), .CK(clock), .Q(SyncY[22]) );
  DFF_X1 \SyncY_reg[21]  ( .D(ElementY[21]), .CK(clock), .Q(SyncY[21]) );
  DFF_X1 \SyncY_reg[20]  ( .D(ElementY[20]), .CK(clock), .Q(SyncY[20]) );
  DFF_X1 \SyncY_reg[19]  ( .D(ElementY[19]), .CK(clock), .Q(SyncY[19]) );
  DFF_X1 \SyncY_reg[18]  ( .D(ElementY[18]), .CK(clock), .Q(SyncY[18]) );
  DFF_X1 \SyncY_reg[17]  ( .D(ElementY[17]), .CK(clock), .Q(SyncY[17]) );
  DFF_X1 \SyncY_reg[16]  ( .D(ElementY[16]), .CK(clock), .Q(SyncY[16]) );
  DFF_X1 \SyncY_reg[15]  ( .D(ElementY[15]), .CK(clock), .Q(SyncY[15]) );
  DFF_X1 \SyncY_reg[14]  ( .D(ElementY[14]), .CK(clock), .Q(SyncY[14]) );
  DFF_X1 \SyncY_reg[13]  ( .D(ElementY[13]), .CK(clock), .Q(SyncY[13]) );
  DFF_X1 \SyncY_reg[12]  ( .D(ElementY[12]), .CK(clock), .Q(SyncY[12]) );
  DFF_X1 \SyncY_reg[11]  ( .D(ElementY[11]), .CK(clock), .Q(SyncY[11]) );
  DFF_X1 \SyncY_reg[10]  ( .D(ElementY[10]), .CK(clock), .Q(SyncY[10]) );
  DFF_X1 \SyncY_reg[9]  ( .D(ElementY[9]), .CK(clock), .Q(SyncY[9]) );
  DFF_X1 \SyncY_reg[8]  ( .D(ElementY[8]), .CK(clock), .Q(SyncY[8]) );
  DFF_X1 \SyncY_reg[7]  ( .D(ElementY[7]), .CK(clock), .Q(SyncY[7]) );
  DFF_X1 \SyncY_reg[6]  ( .D(ElementY[6]), .CK(clock), .Q(SyncY[6]) );
  DFF_X1 \SyncY_reg[5]  ( .D(ElementY[5]), .CK(clock), .Q(SyncY[5]) );
  DFF_X1 \SyncY_reg[4]  ( .D(ElementY[4]), .CK(clock), .Q(SyncY[4]) );
  DFF_X1 \SyncY_reg[3]  ( .D(ElementY[3]), .CK(clock), .Q(SyncY[3]) );
  DFF_X1 \SyncY_reg[2]  ( .D(ElementY[2]), .CK(clock), .Q(SyncY[2]) );
  DFF_X1 \SyncY_reg[1]  ( .D(ElementY[1]), .CK(clock), .Q(SyncY[1]) );
  DFF_X1 \SyncY_reg[0]  ( .D(ElementY[0]), .CK(clock), .Q(SyncY[0]) );
  DFF_X2 \SyncV_reg[0]  ( .D(ElementV[0]), .CK(clock), .Q(SyncV[0]) );
  DFF_X2 \SyncV_reg[1]  ( .D(ElementV[1]), .CK(clock), .Q(SyncV[1]) );
  DFF_X2 \SyncV_reg[2]  ( .D(ElementV[2]), .CK(clock), .Q(SyncV[2]) );
  DFF_X2 \SyncV_reg[3]  ( .D(ElementV[3]), .CK(clock), .Q(SyncV[3]) );
  DFF_X2 \SyncV_reg[4]  ( .D(ElementV[4]), .CK(clock), .Q(SyncV[4]) );
  DFF_X2 \SyncV_reg[5]  ( .D(ElementV[5]), .CK(clock), .Q(SyncV[5]) );
  DFF_X2 \SyncV_reg[6]  ( .D(ElementV[6]), .CK(clock), .Q(SyncV[6]) );
  DFF_X2 \SyncV_reg[7]  ( .D(ElementV[7]), .CK(clock), .Q(SyncV[7]) );
  DFF_X2 \SyncV_reg[8]  ( .D(ElementV[8]), .CK(clock), .Q(SyncV[8]) );
  DFF_X2 \SyncV_reg[9]  ( .D(ElementV[9]), .CK(clock), .Q(SyncV[9]) );
  DFF_X2 \SyncV_reg[10]  ( .D(ElementV[10]), .CK(clock), .Q(SyncV[10]) );
  DFF_X2 \SyncV_reg[11]  ( .D(ElementV[11]), .CK(clock), .Q(SyncV[11]) );
  DFF_X2 \SyncV_reg[12]  ( .D(ElementV[12]), .CK(clock), .Q(SyncV[12]) );
  DFF_X2 \SyncV_reg[13]  ( .D(ElementV[13]), .CK(clock), .Q(SyncV[13]) );
  DFF_X2 \SyncV_reg[14]  ( .D(ElementV[14]), .CK(clock), .Q(SyncV[14]) );
  DFF_X2 \SyncV_reg[15]  ( .D(ElementV[15]), .CK(clock), .Q(SyncV[15]) );
  DFF_X2 \SyncV_reg[16]  ( .D(ElementV[16]), .CK(clock), .Q(SyncV[16]) );
  DFF_X2 \SyncV_reg[17]  ( .D(ElementV[17]), .CK(clock), .Q(SyncV[17]) );
  DFF_X2 \SyncV_reg[18]  ( .D(ElementV[18]), .CK(clock), .Q(SyncV[18]) );
  DFF_X2 \SyncV_reg[19]  ( .D(ElementV[19]), .CK(clock), .Q(SyncV[19]) );
  DFF_X2 \SyncV_reg[20]  ( .D(ElementV[20]), .CK(clock), .Q(SyncV[20]) );
  DFF_X2 \SyncV_reg[21]  ( .D(ElementV[21]), .CK(clock), .Q(SyncV[21]) );
  DFF_X2 \SyncV_reg[22]  ( .D(ElementV[22]), .CK(clock), .Q(SyncV[22]) );
  DFF_X2 \SyncV_reg[23]  ( .D(ElementV[23]), .CK(clock), .Q(SyncV[23]) );
  DFF_X2 \SyncV_reg[24]  ( .D(ElementV[24]), .CK(clock), .Q(SyncV[24]) );
  DFF_X2 \SyncV_reg[25]  ( .D(ElementV[25]), .CK(clock), .Q(SyncV[25]) );
  DFF_X2 \SyncV_reg[26]  ( .D(ElementV[26]), .CK(clock), .Q(SyncV[26]) );
  DFF_X2 \SyncV_reg[27]  ( .D(ElementV[27]), .CK(clock), .Q(SyncV[27]) );
  DFF_X2 \SyncV_reg[28]  ( .D(ElementV[28]), .CK(clock), .Q(SyncV[28]) );
  DFF_X2 \SyncV_reg[29]  ( .D(ElementV[29]), .CK(clock), .Q(SyncV[29]) );
  DFF_X2 \SyncV_reg[30]  ( .D(ElementV[30]), .CK(clock), .Q(SyncV[30]) );
  DFF_X2 \SyncV_reg[31]  ( .D(ElementV[31]), .CK(clock), .Q(SyncV[31]) );
  DFF_X2 \SyncV_reg[32]  ( .D(ElementV[32]), .CK(clock), .Q(SyncV[32]) );
  DFF_X2 \SyncV_reg[33]  ( .D(ElementV[33]), .CK(clock), .Q(SyncV[33]) );
  DFF_X2 \SyncV_reg[34]  ( .D(ElementV[34]), .CK(clock), .Q(SyncV[34]) );
  DFF_X2 \SyncV_reg[35]  ( .D(ElementV[35]), .CK(clock), .Q(SyncV[35]) );
  DFF_X2 \SyncV_reg[36]  ( .D(ElementV[36]), .CK(clock), .Q(SyncV[36]) );
  DFF_X2 \SyncV_reg[37]  ( .D(ElementV[37]), .CK(clock), .Q(SyncV[37]) );
  DFF_X2 \SyncV_reg[38]  ( .D(ElementV[38]), .CK(clock), .Q(SyncV[38]) );
  DFF_X2 \SyncV_reg[39]  ( .D(ElementV[39]), .CK(clock), .Q(SyncV[39]) );
  DFF_X2 \SyncV_reg[40]  ( .D(ElementV[40]), .CK(clock), .Q(SyncV[40]) );
  DFF_X2 \SyncV_reg[41]  ( .D(ElementV[41]), .CK(clock), .Q(SyncV[41]) );
  DFF_X2 \SyncV_reg[42]  ( .D(ElementV[42]), .CK(clock), .Q(SyncV[42]) );
  DFF_X2 \SyncV_reg[43]  ( .D(ElementV[43]), .CK(clock), .Q(SyncV[43]) );
  DFF_X2 \SyncV_reg[44]  ( .D(ElementV[44]), .CK(clock), .Q(SyncV[44]) );
  DFF_X2 \SyncV_reg[45]  ( .D(ElementV[45]), .CK(clock), .Q(SyncV[45]) );
  DFF_X2 \SyncV_reg[46]  ( .D(ElementV[46]), .CK(clock), .Q(SyncV[46]) );
  DFF_X2 \SyncV_reg[47]  ( .D(ElementV[47]), .CK(clock), .Q(SyncV[47]) );
endmodule


module syncDiv ( element1, op1, op2, clock );
  input [47:0] element1;
  output [23:0] op1;
  output [23:0] op2;
  input clock;

  wire   [47:0] buf1;
  wire   [47:0] buf2;
  wire   [47:0] buf3;
  wire   [47:0] buf4;
  wire   [47:0] buf5;
  wire   [47:0] buf6;
  wire   [47:0] buf7;
  wire   [47:0] buf8;
  wire   [47:0] buf9;

  DFF_X1 \buf1_reg[47]  ( .D(element1[47]), .CK(clock), .Q(buf1[47]) );
  DFF_X1 \buf2_reg[47]  ( .D(buf1[47]), .CK(clock), .Q(buf2[47]) );
  DFF_X1 \buf3_reg[47]  ( .D(buf2[47]), .CK(clock), .Q(buf3[47]) );
  DFF_X1 \buf4_reg[47]  ( .D(buf3[47]), .CK(clock), .Q(buf4[47]) );
  DFF_X1 \buf5_reg[47]  ( .D(buf4[47]), .CK(clock), .Q(buf5[47]) );
  DFF_X1 \buf6_reg[47]  ( .D(buf5[47]), .CK(clock), .Q(buf6[47]) );
  DFF_X1 \buf7_reg[47]  ( .D(buf6[47]), .CK(clock), .Q(buf7[47]) );
  DFF_X1 \buf8_reg[47]  ( .D(buf7[47]), .CK(clock), .Q(buf8[47]) );
  DFF_X1 \buf9_reg[47]  ( .D(buf8[47]), .CK(clock), .Q(buf9[47]) );
  DFF_X1 \buf1_reg[46]  ( .D(element1[46]), .CK(clock), .Q(buf1[46]) );
  DFF_X1 \buf2_reg[46]  ( .D(buf1[46]), .CK(clock), .Q(buf2[46]) );
  DFF_X1 \buf3_reg[46]  ( .D(buf2[46]), .CK(clock), .Q(buf3[46]) );
  DFF_X1 \buf4_reg[46]  ( .D(buf3[46]), .CK(clock), .Q(buf4[46]) );
  DFF_X1 \buf5_reg[46]  ( .D(buf4[46]), .CK(clock), .Q(buf5[46]) );
  DFF_X1 \buf6_reg[46]  ( .D(buf5[46]), .CK(clock), .Q(buf6[46]) );
  DFF_X1 \buf7_reg[46]  ( .D(buf6[46]), .CK(clock), .Q(buf7[46]) );
  DFF_X1 \buf8_reg[46]  ( .D(buf7[46]), .CK(clock), .Q(buf8[46]) );
  DFF_X1 \buf9_reg[46]  ( .D(buf8[46]), .CK(clock), .Q(buf9[46]) );
  DFF_X1 \buf1_reg[45]  ( .D(element1[45]), .CK(clock), .Q(buf1[45]) );
  DFF_X1 \buf2_reg[45]  ( .D(buf1[45]), .CK(clock), .Q(buf2[45]) );
  DFF_X1 \buf3_reg[45]  ( .D(buf2[45]), .CK(clock), .Q(buf3[45]) );
  DFF_X1 \buf4_reg[45]  ( .D(buf3[45]), .CK(clock), .Q(buf4[45]) );
  DFF_X1 \buf5_reg[45]  ( .D(buf4[45]), .CK(clock), .Q(buf5[45]) );
  DFF_X1 \buf6_reg[45]  ( .D(buf5[45]), .CK(clock), .Q(buf6[45]) );
  DFF_X1 \buf7_reg[45]  ( .D(buf6[45]), .CK(clock), .Q(buf7[45]) );
  DFF_X1 \buf8_reg[45]  ( .D(buf7[45]), .CK(clock), .Q(buf8[45]) );
  DFF_X1 \buf9_reg[45]  ( .D(buf8[45]), .CK(clock), .Q(buf9[45]) );
  DFF_X1 \buf1_reg[44]  ( .D(element1[44]), .CK(clock), .Q(buf1[44]) );
  DFF_X1 \buf2_reg[44]  ( .D(buf1[44]), .CK(clock), .Q(buf2[44]) );
  DFF_X1 \buf3_reg[44]  ( .D(buf2[44]), .CK(clock), .Q(buf3[44]) );
  DFF_X1 \buf4_reg[44]  ( .D(buf3[44]), .CK(clock), .Q(buf4[44]) );
  DFF_X1 \buf5_reg[44]  ( .D(buf4[44]), .CK(clock), .Q(buf5[44]) );
  DFF_X1 \buf6_reg[44]  ( .D(buf5[44]), .CK(clock), .Q(buf6[44]) );
  DFF_X1 \buf7_reg[44]  ( .D(buf6[44]), .CK(clock), .Q(buf7[44]) );
  DFF_X1 \buf8_reg[44]  ( .D(buf7[44]), .CK(clock), .Q(buf8[44]) );
  DFF_X1 \buf9_reg[44]  ( .D(buf8[44]), .CK(clock), .Q(buf9[44]) );
  DFF_X1 \buf1_reg[43]  ( .D(element1[43]), .CK(clock), .Q(buf1[43]) );
  DFF_X1 \buf2_reg[43]  ( .D(buf1[43]), .CK(clock), .Q(buf2[43]) );
  DFF_X1 \buf3_reg[43]  ( .D(buf2[43]), .CK(clock), .Q(buf3[43]) );
  DFF_X1 \buf4_reg[43]  ( .D(buf3[43]), .CK(clock), .Q(buf4[43]) );
  DFF_X1 \buf5_reg[43]  ( .D(buf4[43]), .CK(clock), .Q(buf5[43]) );
  DFF_X1 \buf6_reg[43]  ( .D(buf5[43]), .CK(clock), .Q(buf6[43]) );
  DFF_X1 \buf7_reg[43]  ( .D(buf6[43]), .CK(clock), .Q(buf7[43]) );
  DFF_X1 \buf8_reg[43]  ( .D(buf7[43]), .CK(clock), .Q(buf8[43]) );
  DFF_X1 \buf9_reg[43]  ( .D(buf8[43]), .CK(clock), .Q(buf9[43]) );
  DFF_X1 \buf1_reg[42]  ( .D(element1[42]), .CK(clock), .Q(buf1[42]) );
  DFF_X1 \buf2_reg[42]  ( .D(buf1[42]), .CK(clock), .Q(buf2[42]) );
  DFF_X1 \buf3_reg[42]  ( .D(buf2[42]), .CK(clock), .Q(buf3[42]) );
  DFF_X1 \buf4_reg[42]  ( .D(buf3[42]), .CK(clock), .Q(buf4[42]) );
  DFF_X1 \buf5_reg[42]  ( .D(buf4[42]), .CK(clock), .Q(buf5[42]) );
  DFF_X1 \buf6_reg[42]  ( .D(buf5[42]), .CK(clock), .Q(buf6[42]) );
  DFF_X1 \buf7_reg[42]  ( .D(buf6[42]), .CK(clock), .Q(buf7[42]) );
  DFF_X1 \buf8_reg[42]  ( .D(buf7[42]), .CK(clock), .Q(buf8[42]) );
  DFF_X1 \buf9_reg[42]  ( .D(buf8[42]), .CK(clock), .Q(buf9[42]) );
  DFF_X1 \buf1_reg[41]  ( .D(element1[41]), .CK(clock), .Q(buf1[41]) );
  DFF_X1 \buf2_reg[41]  ( .D(buf1[41]), .CK(clock), .Q(buf2[41]) );
  DFF_X1 \buf3_reg[41]  ( .D(buf2[41]), .CK(clock), .Q(buf3[41]) );
  DFF_X1 \buf4_reg[41]  ( .D(buf3[41]), .CK(clock), .Q(buf4[41]) );
  DFF_X1 \buf5_reg[41]  ( .D(buf4[41]), .CK(clock), .Q(buf5[41]) );
  DFF_X1 \buf6_reg[41]  ( .D(buf5[41]), .CK(clock), .Q(buf6[41]) );
  DFF_X1 \buf7_reg[41]  ( .D(buf6[41]), .CK(clock), .Q(buf7[41]) );
  DFF_X1 \buf8_reg[41]  ( .D(buf7[41]), .CK(clock), .Q(buf8[41]) );
  DFF_X1 \buf9_reg[41]  ( .D(buf8[41]), .CK(clock), .Q(buf9[41]) );
  DFF_X1 \buf1_reg[40]  ( .D(element1[40]), .CK(clock), .Q(buf1[40]) );
  DFF_X1 \buf2_reg[40]  ( .D(buf1[40]), .CK(clock), .Q(buf2[40]) );
  DFF_X1 \buf3_reg[40]  ( .D(buf2[40]), .CK(clock), .Q(buf3[40]) );
  DFF_X1 \buf4_reg[40]  ( .D(buf3[40]), .CK(clock), .Q(buf4[40]) );
  DFF_X1 \buf5_reg[40]  ( .D(buf4[40]), .CK(clock), .Q(buf5[40]) );
  DFF_X1 \buf6_reg[40]  ( .D(buf5[40]), .CK(clock), .Q(buf6[40]) );
  DFF_X1 \buf7_reg[40]  ( .D(buf6[40]), .CK(clock), .Q(buf7[40]) );
  DFF_X1 \buf8_reg[40]  ( .D(buf7[40]), .CK(clock), .Q(buf8[40]) );
  DFF_X1 \buf9_reg[40]  ( .D(buf8[40]), .CK(clock), .Q(buf9[40]) );
  DFF_X1 \buf1_reg[39]  ( .D(element1[39]), .CK(clock), .Q(buf1[39]) );
  DFF_X1 \buf2_reg[39]  ( .D(buf1[39]), .CK(clock), .Q(buf2[39]) );
  DFF_X1 \buf3_reg[39]  ( .D(buf2[39]), .CK(clock), .Q(buf3[39]) );
  DFF_X1 \buf4_reg[39]  ( .D(buf3[39]), .CK(clock), .Q(buf4[39]) );
  DFF_X1 \buf5_reg[39]  ( .D(buf4[39]), .CK(clock), .Q(buf5[39]) );
  DFF_X1 \buf6_reg[39]  ( .D(buf5[39]), .CK(clock), .Q(buf6[39]) );
  DFF_X1 \buf7_reg[39]  ( .D(buf6[39]), .CK(clock), .Q(buf7[39]) );
  DFF_X1 \buf8_reg[39]  ( .D(buf7[39]), .CK(clock), .Q(buf8[39]) );
  DFF_X1 \buf9_reg[39]  ( .D(buf8[39]), .CK(clock), .Q(buf9[39]) );
  DFF_X1 \buf1_reg[38]  ( .D(element1[38]), .CK(clock), .Q(buf1[38]) );
  DFF_X1 \buf2_reg[38]  ( .D(buf1[38]), .CK(clock), .Q(buf2[38]) );
  DFF_X1 \buf3_reg[38]  ( .D(buf2[38]), .CK(clock), .Q(buf3[38]) );
  DFF_X1 \buf4_reg[38]  ( .D(buf3[38]), .CK(clock), .Q(buf4[38]) );
  DFF_X1 \buf5_reg[38]  ( .D(buf4[38]), .CK(clock), .Q(buf5[38]) );
  DFF_X1 \buf6_reg[38]  ( .D(buf5[38]), .CK(clock), .Q(buf6[38]) );
  DFF_X1 \buf7_reg[38]  ( .D(buf6[38]), .CK(clock), .Q(buf7[38]) );
  DFF_X1 \buf8_reg[38]  ( .D(buf7[38]), .CK(clock), .Q(buf8[38]) );
  DFF_X1 \buf9_reg[38]  ( .D(buf8[38]), .CK(clock), .Q(buf9[38]) );
  DFF_X1 \buf1_reg[37]  ( .D(element1[37]), .CK(clock), .Q(buf1[37]) );
  DFF_X1 \buf2_reg[37]  ( .D(buf1[37]), .CK(clock), .Q(buf2[37]) );
  DFF_X1 \buf3_reg[37]  ( .D(buf2[37]), .CK(clock), .Q(buf3[37]) );
  DFF_X1 \buf4_reg[37]  ( .D(buf3[37]), .CK(clock), .Q(buf4[37]) );
  DFF_X1 \buf5_reg[37]  ( .D(buf4[37]), .CK(clock), .Q(buf5[37]) );
  DFF_X1 \buf6_reg[37]  ( .D(buf5[37]), .CK(clock), .Q(buf6[37]) );
  DFF_X1 \buf7_reg[37]  ( .D(buf6[37]), .CK(clock), .Q(buf7[37]) );
  DFF_X1 \buf8_reg[37]  ( .D(buf7[37]), .CK(clock), .Q(buf8[37]) );
  DFF_X1 \buf9_reg[37]  ( .D(buf8[37]), .CK(clock), .Q(buf9[37]) );
  DFF_X1 \buf1_reg[36]  ( .D(element1[36]), .CK(clock), .Q(buf1[36]) );
  DFF_X1 \buf2_reg[36]  ( .D(buf1[36]), .CK(clock), .Q(buf2[36]) );
  DFF_X1 \buf3_reg[36]  ( .D(buf2[36]), .CK(clock), .Q(buf3[36]) );
  DFF_X1 \buf4_reg[36]  ( .D(buf3[36]), .CK(clock), .Q(buf4[36]) );
  DFF_X1 \buf5_reg[36]  ( .D(buf4[36]), .CK(clock), .Q(buf5[36]) );
  DFF_X1 \buf6_reg[36]  ( .D(buf5[36]), .CK(clock), .Q(buf6[36]) );
  DFF_X1 \buf7_reg[36]  ( .D(buf6[36]), .CK(clock), .Q(buf7[36]) );
  DFF_X1 \buf8_reg[36]  ( .D(buf7[36]), .CK(clock), .Q(buf8[36]) );
  DFF_X1 \buf9_reg[36]  ( .D(buf8[36]), .CK(clock), .Q(buf9[36]) );
  DFF_X1 \buf1_reg[35]  ( .D(element1[35]), .CK(clock), .Q(buf1[35]) );
  DFF_X1 \buf2_reg[35]  ( .D(buf1[35]), .CK(clock), .Q(buf2[35]) );
  DFF_X1 \buf3_reg[35]  ( .D(buf2[35]), .CK(clock), .Q(buf3[35]) );
  DFF_X1 \buf4_reg[35]  ( .D(buf3[35]), .CK(clock), .Q(buf4[35]) );
  DFF_X1 \buf5_reg[35]  ( .D(buf4[35]), .CK(clock), .Q(buf5[35]) );
  DFF_X1 \buf6_reg[35]  ( .D(buf5[35]), .CK(clock), .Q(buf6[35]) );
  DFF_X1 \buf7_reg[35]  ( .D(buf6[35]), .CK(clock), .Q(buf7[35]) );
  DFF_X1 \buf8_reg[35]  ( .D(buf7[35]), .CK(clock), .Q(buf8[35]) );
  DFF_X1 \buf9_reg[35]  ( .D(buf8[35]), .CK(clock), .Q(buf9[35]) );
  DFF_X1 \buf1_reg[34]  ( .D(element1[34]), .CK(clock), .Q(buf1[34]) );
  DFF_X1 \buf2_reg[34]  ( .D(buf1[34]), .CK(clock), .Q(buf2[34]) );
  DFF_X1 \buf3_reg[34]  ( .D(buf2[34]), .CK(clock), .Q(buf3[34]) );
  DFF_X1 \buf4_reg[34]  ( .D(buf3[34]), .CK(clock), .Q(buf4[34]) );
  DFF_X1 \buf5_reg[34]  ( .D(buf4[34]), .CK(clock), .Q(buf5[34]) );
  DFF_X1 \buf6_reg[34]  ( .D(buf5[34]), .CK(clock), .Q(buf6[34]) );
  DFF_X1 \buf7_reg[34]  ( .D(buf6[34]), .CK(clock), .Q(buf7[34]) );
  DFF_X1 \buf8_reg[34]  ( .D(buf7[34]), .CK(clock), .Q(buf8[34]) );
  DFF_X1 \buf9_reg[34]  ( .D(buf8[34]), .CK(clock), .Q(buf9[34]) );
  DFF_X1 \buf1_reg[33]  ( .D(element1[33]), .CK(clock), .Q(buf1[33]) );
  DFF_X1 \buf2_reg[33]  ( .D(buf1[33]), .CK(clock), .Q(buf2[33]) );
  DFF_X1 \buf3_reg[33]  ( .D(buf2[33]), .CK(clock), .Q(buf3[33]) );
  DFF_X1 \buf4_reg[33]  ( .D(buf3[33]), .CK(clock), .Q(buf4[33]) );
  DFF_X1 \buf5_reg[33]  ( .D(buf4[33]), .CK(clock), .Q(buf5[33]) );
  DFF_X1 \buf6_reg[33]  ( .D(buf5[33]), .CK(clock), .Q(buf6[33]) );
  DFF_X1 \buf7_reg[33]  ( .D(buf6[33]), .CK(clock), .Q(buf7[33]) );
  DFF_X1 \buf8_reg[33]  ( .D(buf7[33]), .CK(clock), .Q(buf8[33]) );
  DFF_X1 \buf9_reg[33]  ( .D(buf8[33]), .CK(clock), .Q(buf9[33]) );
  DFF_X1 \buf1_reg[32]  ( .D(element1[32]), .CK(clock), .Q(buf1[32]) );
  DFF_X1 \buf2_reg[32]  ( .D(buf1[32]), .CK(clock), .Q(buf2[32]) );
  DFF_X1 \buf3_reg[32]  ( .D(buf2[32]), .CK(clock), .Q(buf3[32]) );
  DFF_X1 \buf4_reg[32]  ( .D(buf3[32]), .CK(clock), .Q(buf4[32]) );
  DFF_X1 \buf5_reg[32]  ( .D(buf4[32]), .CK(clock), .Q(buf5[32]) );
  DFF_X1 \buf6_reg[32]  ( .D(buf5[32]), .CK(clock), .Q(buf6[32]) );
  DFF_X1 \buf7_reg[32]  ( .D(buf6[32]), .CK(clock), .Q(buf7[32]) );
  DFF_X1 \buf8_reg[32]  ( .D(buf7[32]), .CK(clock), .Q(buf8[32]) );
  DFF_X1 \buf9_reg[32]  ( .D(buf8[32]), .CK(clock), .Q(buf9[32]) );
  DFF_X1 \buf1_reg[31]  ( .D(element1[31]), .CK(clock), .Q(buf1[31]) );
  DFF_X1 \buf2_reg[31]  ( .D(buf1[31]), .CK(clock), .Q(buf2[31]) );
  DFF_X1 \buf3_reg[31]  ( .D(buf2[31]), .CK(clock), .Q(buf3[31]) );
  DFF_X1 \buf4_reg[31]  ( .D(buf3[31]), .CK(clock), .Q(buf4[31]) );
  DFF_X1 \buf5_reg[31]  ( .D(buf4[31]), .CK(clock), .Q(buf5[31]) );
  DFF_X1 \buf6_reg[31]  ( .D(buf5[31]), .CK(clock), .Q(buf6[31]) );
  DFF_X1 \buf7_reg[31]  ( .D(buf6[31]), .CK(clock), .Q(buf7[31]) );
  DFF_X1 \buf8_reg[31]  ( .D(buf7[31]), .CK(clock), .Q(buf8[31]) );
  DFF_X1 \buf9_reg[31]  ( .D(buf8[31]), .CK(clock), .Q(buf9[31]) );
  DFF_X1 \buf1_reg[30]  ( .D(element1[30]), .CK(clock), .Q(buf1[30]) );
  DFF_X1 \buf2_reg[30]  ( .D(buf1[30]), .CK(clock), .Q(buf2[30]) );
  DFF_X1 \buf3_reg[30]  ( .D(buf2[30]), .CK(clock), .Q(buf3[30]) );
  DFF_X1 \buf4_reg[30]  ( .D(buf3[30]), .CK(clock), .Q(buf4[30]) );
  DFF_X1 \buf5_reg[30]  ( .D(buf4[30]), .CK(clock), .Q(buf5[30]) );
  DFF_X1 \buf6_reg[30]  ( .D(buf5[30]), .CK(clock), .Q(buf6[30]) );
  DFF_X1 \buf7_reg[30]  ( .D(buf6[30]), .CK(clock), .Q(buf7[30]) );
  DFF_X1 \buf8_reg[30]  ( .D(buf7[30]), .CK(clock), .Q(buf8[30]) );
  DFF_X1 \buf9_reg[30]  ( .D(buf8[30]), .CK(clock), .Q(buf9[30]) );
  DFF_X1 \buf1_reg[29]  ( .D(element1[29]), .CK(clock), .Q(buf1[29]) );
  DFF_X1 \buf2_reg[29]  ( .D(buf1[29]), .CK(clock), .Q(buf2[29]) );
  DFF_X1 \buf3_reg[29]  ( .D(buf2[29]), .CK(clock), .Q(buf3[29]) );
  DFF_X1 \buf4_reg[29]  ( .D(buf3[29]), .CK(clock), .Q(buf4[29]) );
  DFF_X1 \buf5_reg[29]  ( .D(buf4[29]), .CK(clock), .Q(buf5[29]) );
  DFF_X1 \buf6_reg[29]  ( .D(buf5[29]), .CK(clock), .Q(buf6[29]) );
  DFF_X1 \buf7_reg[29]  ( .D(buf6[29]), .CK(clock), .Q(buf7[29]) );
  DFF_X1 \buf8_reg[29]  ( .D(buf7[29]), .CK(clock), .Q(buf8[29]) );
  DFF_X1 \buf9_reg[29]  ( .D(buf8[29]), .CK(clock), .Q(buf9[29]) );
  DFF_X1 \buf1_reg[28]  ( .D(element1[28]), .CK(clock), .Q(buf1[28]) );
  DFF_X1 \buf2_reg[28]  ( .D(buf1[28]), .CK(clock), .Q(buf2[28]) );
  DFF_X1 \buf3_reg[28]  ( .D(buf2[28]), .CK(clock), .Q(buf3[28]) );
  DFF_X1 \buf4_reg[28]  ( .D(buf3[28]), .CK(clock), .Q(buf4[28]) );
  DFF_X1 \buf5_reg[28]  ( .D(buf4[28]), .CK(clock), .Q(buf5[28]) );
  DFF_X1 \buf6_reg[28]  ( .D(buf5[28]), .CK(clock), .Q(buf6[28]) );
  DFF_X1 \buf7_reg[28]  ( .D(buf6[28]), .CK(clock), .Q(buf7[28]) );
  DFF_X1 \buf8_reg[28]  ( .D(buf7[28]), .CK(clock), .Q(buf8[28]) );
  DFF_X1 \buf9_reg[28]  ( .D(buf8[28]), .CK(clock), .Q(buf9[28]) );
  DFF_X1 \buf1_reg[27]  ( .D(element1[27]), .CK(clock), .Q(buf1[27]) );
  DFF_X1 \buf2_reg[27]  ( .D(buf1[27]), .CK(clock), .Q(buf2[27]) );
  DFF_X1 \buf3_reg[27]  ( .D(buf2[27]), .CK(clock), .Q(buf3[27]) );
  DFF_X1 \buf4_reg[27]  ( .D(buf3[27]), .CK(clock), .Q(buf4[27]) );
  DFF_X1 \buf5_reg[27]  ( .D(buf4[27]), .CK(clock), .Q(buf5[27]) );
  DFF_X1 \buf6_reg[27]  ( .D(buf5[27]), .CK(clock), .Q(buf6[27]) );
  DFF_X1 \buf7_reg[27]  ( .D(buf6[27]), .CK(clock), .Q(buf7[27]) );
  DFF_X1 \buf8_reg[27]  ( .D(buf7[27]), .CK(clock), .Q(buf8[27]) );
  DFF_X1 \buf9_reg[27]  ( .D(buf8[27]), .CK(clock), .Q(buf9[27]) );
  DFF_X1 \buf1_reg[26]  ( .D(element1[26]), .CK(clock), .Q(buf1[26]) );
  DFF_X1 \buf2_reg[26]  ( .D(buf1[26]), .CK(clock), .Q(buf2[26]) );
  DFF_X1 \buf3_reg[26]  ( .D(buf2[26]), .CK(clock), .Q(buf3[26]) );
  DFF_X1 \buf4_reg[26]  ( .D(buf3[26]), .CK(clock), .Q(buf4[26]) );
  DFF_X1 \buf5_reg[26]  ( .D(buf4[26]), .CK(clock), .Q(buf5[26]) );
  DFF_X1 \buf6_reg[26]  ( .D(buf5[26]), .CK(clock), .Q(buf6[26]) );
  DFF_X1 \buf7_reg[26]  ( .D(buf6[26]), .CK(clock), .Q(buf7[26]) );
  DFF_X1 \buf8_reg[26]  ( .D(buf7[26]), .CK(clock), .Q(buf8[26]) );
  DFF_X1 \buf9_reg[26]  ( .D(buf8[26]), .CK(clock), .Q(buf9[26]) );
  DFF_X1 \buf1_reg[25]  ( .D(element1[25]), .CK(clock), .Q(buf1[25]) );
  DFF_X1 \buf2_reg[25]  ( .D(buf1[25]), .CK(clock), .Q(buf2[25]) );
  DFF_X1 \buf3_reg[25]  ( .D(buf2[25]), .CK(clock), .Q(buf3[25]) );
  DFF_X1 \buf4_reg[25]  ( .D(buf3[25]), .CK(clock), .Q(buf4[25]) );
  DFF_X1 \buf5_reg[25]  ( .D(buf4[25]), .CK(clock), .Q(buf5[25]) );
  DFF_X1 \buf6_reg[25]  ( .D(buf5[25]), .CK(clock), .Q(buf6[25]) );
  DFF_X1 \buf7_reg[25]  ( .D(buf6[25]), .CK(clock), .Q(buf7[25]) );
  DFF_X1 \buf8_reg[25]  ( .D(buf7[25]), .CK(clock), .Q(buf8[25]) );
  DFF_X1 \buf9_reg[25]  ( .D(buf8[25]), .CK(clock), .Q(buf9[25]) );
  DFF_X1 \buf1_reg[24]  ( .D(element1[24]), .CK(clock), .Q(buf1[24]) );
  DFF_X1 \buf2_reg[24]  ( .D(buf1[24]), .CK(clock), .Q(buf2[24]) );
  DFF_X1 \buf3_reg[24]  ( .D(buf2[24]), .CK(clock), .Q(buf3[24]) );
  DFF_X1 \buf4_reg[24]  ( .D(buf3[24]), .CK(clock), .Q(buf4[24]) );
  DFF_X1 \buf5_reg[24]  ( .D(buf4[24]), .CK(clock), .Q(buf5[24]) );
  DFF_X1 \buf6_reg[24]  ( .D(buf5[24]), .CK(clock), .Q(buf6[24]) );
  DFF_X1 \buf7_reg[24]  ( .D(buf6[24]), .CK(clock), .Q(buf7[24]) );
  DFF_X1 \buf8_reg[24]  ( .D(buf7[24]), .CK(clock), .Q(buf8[24]) );
  DFF_X1 \buf9_reg[24]  ( .D(buf8[24]), .CK(clock), .Q(buf9[24]) );
  DFF_X1 \buf1_reg[23]  ( .D(element1[23]), .CK(clock), .Q(buf1[23]) );
  DFF_X1 \buf2_reg[23]  ( .D(buf1[23]), .CK(clock), .Q(buf2[23]) );
  DFF_X1 \buf3_reg[23]  ( .D(buf2[23]), .CK(clock), .Q(buf3[23]) );
  DFF_X1 \buf4_reg[23]  ( .D(buf3[23]), .CK(clock), .Q(buf4[23]) );
  DFF_X1 \buf5_reg[23]  ( .D(buf4[23]), .CK(clock), .Q(buf5[23]) );
  DFF_X1 \buf6_reg[23]  ( .D(buf5[23]), .CK(clock), .Q(buf6[23]) );
  DFF_X1 \buf7_reg[23]  ( .D(buf6[23]), .CK(clock), .Q(buf7[23]) );
  DFF_X1 \buf8_reg[23]  ( .D(buf7[23]), .CK(clock), .Q(buf8[23]) );
  DFF_X1 \buf9_reg[23]  ( .D(buf8[23]), .CK(clock), .Q(buf9[23]) );
  DFF_X1 \buf1_reg[22]  ( .D(element1[22]), .CK(clock), .Q(buf1[22]) );
  DFF_X1 \buf2_reg[22]  ( .D(buf1[22]), .CK(clock), .Q(buf2[22]) );
  DFF_X1 \buf3_reg[22]  ( .D(buf2[22]), .CK(clock), .Q(buf3[22]) );
  DFF_X1 \buf4_reg[22]  ( .D(buf3[22]), .CK(clock), .Q(buf4[22]) );
  DFF_X1 \buf5_reg[22]  ( .D(buf4[22]), .CK(clock), .Q(buf5[22]) );
  DFF_X1 \buf6_reg[22]  ( .D(buf5[22]), .CK(clock), .Q(buf6[22]) );
  DFF_X1 \buf7_reg[22]  ( .D(buf6[22]), .CK(clock), .Q(buf7[22]) );
  DFF_X1 \buf8_reg[22]  ( .D(buf7[22]), .CK(clock), .Q(buf8[22]) );
  DFF_X1 \buf9_reg[22]  ( .D(buf8[22]), .CK(clock), .Q(buf9[22]) );
  DFF_X1 \buf1_reg[21]  ( .D(element1[21]), .CK(clock), .Q(buf1[21]) );
  DFF_X1 \buf2_reg[21]  ( .D(buf1[21]), .CK(clock), .Q(buf2[21]) );
  DFF_X1 \buf3_reg[21]  ( .D(buf2[21]), .CK(clock), .Q(buf3[21]) );
  DFF_X1 \buf4_reg[21]  ( .D(buf3[21]), .CK(clock), .Q(buf4[21]) );
  DFF_X1 \buf5_reg[21]  ( .D(buf4[21]), .CK(clock), .Q(buf5[21]) );
  DFF_X1 \buf6_reg[21]  ( .D(buf5[21]), .CK(clock), .Q(buf6[21]) );
  DFF_X1 \buf7_reg[21]  ( .D(buf6[21]), .CK(clock), .Q(buf7[21]) );
  DFF_X1 \buf8_reg[21]  ( .D(buf7[21]), .CK(clock), .Q(buf8[21]) );
  DFF_X1 \buf9_reg[21]  ( .D(buf8[21]), .CK(clock), .Q(buf9[21]) );
  DFF_X1 \buf1_reg[20]  ( .D(element1[20]), .CK(clock), .Q(buf1[20]) );
  DFF_X1 \buf2_reg[20]  ( .D(buf1[20]), .CK(clock), .Q(buf2[20]) );
  DFF_X1 \buf3_reg[20]  ( .D(buf2[20]), .CK(clock), .Q(buf3[20]) );
  DFF_X1 \buf4_reg[20]  ( .D(buf3[20]), .CK(clock), .Q(buf4[20]) );
  DFF_X1 \buf5_reg[20]  ( .D(buf4[20]), .CK(clock), .Q(buf5[20]) );
  DFF_X1 \buf6_reg[20]  ( .D(buf5[20]), .CK(clock), .Q(buf6[20]) );
  DFF_X1 \buf7_reg[20]  ( .D(buf6[20]), .CK(clock), .Q(buf7[20]) );
  DFF_X1 \buf8_reg[20]  ( .D(buf7[20]), .CK(clock), .Q(buf8[20]) );
  DFF_X1 \buf9_reg[20]  ( .D(buf8[20]), .CK(clock), .Q(buf9[20]) );
  DFF_X1 \buf1_reg[19]  ( .D(element1[19]), .CK(clock), .Q(buf1[19]) );
  DFF_X1 \buf2_reg[19]  ( .D(buf1[19]), .CK(clock), .Q(buf2[19]) );
  DFF_X1 \buf3_reg[19]  ( .D(buf2[19]), .CK(clock), .Q(buf3[19]) );
  DFF_X1 \buf4_reg[19]  ( .D(buf3[19]), .CK(clock), .Q(buf4[19]) );
  DFF_X1 \buf5_reg[19]  ( .D(buf4[19]), .CK(clock), .Q(buf5[19]) );
  DFF_X1 \buf6_reg[19]  ( .D(buf5[19]), .CK(clock), .Q(buf6[19]) );
  DFF_X1 \buf7_reg[19]  ( .D(buf6[19]), .CK(clock), .Q(buf7[19]) );
  DFF_X1 \buf8_reg[19]  ( .D(buf7[19]), .CK(clock), .Q(buf8[19]) );
  DFF_X1 \buf9_reg[19]  ( .D(buf8[19]), .CK(clock), .Q(buf9[19]) );
  DFF_X1 \buf1_reg[18]  ( .D(element1[18]), .CK(clock), .Q(buf1[18]) );
  DFF_X1 \buf2_reg[18]  ( .D(buf1[18]), .CK(clock), .Q(buf2[18]) );
  DFF_X1 \buf3_reg[18]  ( .D(buf2[18]), .CK(clock), .Q(buf3[18]) );
  DFF_X1 \buf4_reg[18]  ( .D(buf3[18]), .CK(clock), .Q(buf4[18]) );
  DFF_X1 \buf5_reg[18]  ( .D(buf4[18]), .CK(clock), .Q(buf5[18]) );
  DFF_X1 \buf6_reg[18]  ( .D(buf5[18]), .CK(clock), .Q(buf6[18]) );
  DFF_X1 \buf7_reg[18]  ( .D(buf6[18]), .CK(clock), .Q(buf7[18]) );
  DFF_X1 \buf8_reg[18]  ( .D(buf7[18]), .CK(clock), .Q(buf8[18]) );
  DFF_X1 \buf9_reg[18]  ( .D(buf8[18]), .CK(clock), .Q(buf9[18]) );
  DFF_X1 \buf1_reg[17]  ( .D(element1[17]), .CK(clock), .Q(buf1[17]) );
  DFF_X1 \buf2_reg[17]  ( .D(buf1[17]), .CK(clock), .Q(buf2[17]) );
  DFF_X1 \buf3_reg[17]  ( .D(buf2[17]), .CK(clock), .Q(buf3[17]) );
  DFF_X1 \buf4_reg[17]  ( .D(buf3[17]), .CK(clock), .Q(buf4[17]) );
  DFF_X1 \buf5_reg[17]  ( .D(buf4[17]), .CK(clock), .Q(buf5[17]) );
  DFF_X1 \buf6_reg[17]  ( .D(buf5[17]), .CK(clock), .Q(buf6[17]) );
  DFF_X1 \buf7_reg[17]  ( .D(buf6[17]), .CK(clock), .Q(buf7[17]) );
  DFF_X1 \buf8_reg[17]  ( .D(buf7[17]), .CK(clock), .Q(buf8[17]) );
  DFF_X1 \buf9_reg[17]  ( .D(buf8[17]), .CK(clock), .Q(buf9[17]) );
  DFF_X1 \buf1_reg[16]  ( .D(element1[16]), .CK(clock), .Q(buf1[16]) );
  DFF_X1 \buf2_reg[16]  ( .D(buf1[16]), .CK(clock), .Q(buf2[16]) );
  DFF_X1 \buf3_reg[16]  ( .D(buf2[16]), .CK(clock), .Q(buf3[16]) );
  DFF_X1 \buf4_reg[16]  ( .D(buf3[16]), .CK(clock), .Q(buf4[16]) );
  DFF_X1 \buf5_reg[16]  ( .D(buf4[16]), .CK(clock), .Q(buf5[16]) );
  DFF_X1 \buf6_reg[16]  ( .D(buf5[16]), .CK(clock), .Q(buf6[16]) );
  DFF_X1 \buf7_reg[16]  ( .D(buf6[16]), .CK(clock), .Q(buf7[16]) );
  DFF_X1 \buf8_reg[16]  ( .D(buf7[16]), .CK(clock), .Q(buf8[16]) );
  DFF_X1 \buf9_reg[16]  ( .D(buf8[16]), .CK(clock), .Q(buf9[16]) );
  DFF_X1 \buf1_reg[15]  ( .D(element1[15]), .CK(clock), .Q(buf1[15]) );
  DFF_X1 \buf2_reg[15]  ( .D(buf1[15]), .CK(clock), .Q(buf2[15]) );
  DFF_X1 \buf3_reg[15]  ( .D(buf2[15]), .CK(clock), .Q(buf3[15]) );
  DFF_X1 \buf4_reg[15]  ( .D(buf3[15]), .CK(clock), .Q(buf4[15]) );
  DFF_X1 \buf5_reg[15]  ( .D(buf4[15]), .CK(clock), .Q(buf5[15]) );
  DFF_X1 \buf6_reg[15]  ( .D(buf5[15]), .CK(clock), .Q(buf6[15]) );
  DFF_X1 \buf7_reg[15]  ( .D(buf6[15]), .CK(clock), .Q(buf7[15]) );
  DFF_X1 \buf8_reg[15]  ( .D(buf7[15]), .CK(clock), .Q(buf8[15]) );
  DFF_X1 \buf9_reg[15]  ( .D(buf8[15]), .CK(clock), .Q(buf9[15]) );
  DFF_X1 \buf1_reg[14]  ( .D(element1[14]), .CK(clock), .Q(buf1[14]) );
  DFF_X1 \buf2_reg[14]  ( .D(buf1[14]), .CK(clock), .Q(buf2[14]) );
  DFF_X1 \buf3_reg[14]  ( .D(buf2[14]), .CK(clock), .Q(buf3[14]) );
  DFF_X1 \buf4_reg[14]  ( .D(buf3[14]), .CK(clock), .Q(buf4[14]) );
  DFF_X1 \buf5_reg[14]  ( .D(buf4[14]), .CK(clock), .Q(buf5[14]) );
  DFF_X1 \buf6_reg[14]  ( .D(buf5[14]), .CK(clock), .Q(buf6[14]) );
  DFF_X1 \buf7_reg[14]  ( .D(buf6[14]), .CK(clock), .Q(buf7[14]) );
  DFF_X1 \buf8_reg[14]  ( .D(buf7[14]), .CK(clock), .Q(buf8[14]) );
  DFF_X1 \buf9_reg[14]  ( .D(buf8[14]), .CK(clock), .Q(buf9[14]) );
  DFF_X1 \buf1_reg[13]  ( .D(element1[13]), .CK(clock), .Q(buf1[13]) );
  DFF_X1 \buf2_reg[13]  ( .D(buf1[13]), .CK(clock), .Q(buf2[13]) );
  DFF_X1 \buf3_reg[13]  ( .D(buf2[13]), .CK(clock), .Q(buf3[13]) );
  DFF_X1 \buf4_reg[13]  ( .D(buf3[13]), .CK(clock), .Q(buf4[13]) );
  DFF_X1 \buf5_reg[13]  ( .D(buf4[13]), .CK(clock), .Q(buf5[13]) );
  DFF_X1 \buf6_reg[13]  ( .D(buf5[13]), .CK(clock), .Q(buf6[13]) );
  DFF_X1 \buf7_reg[13]  ( .D(buf6[13]), .CK(clock), .Q(buf7[13]) );
  DFF_X1 \buf8_reg[13]  ( .D(buf7[13]), .CK(clock), .Q(buf8[13]) );
  DFF_X1 \buf9_reg[13]  ( .D(buf8[13]), .CK(clock), .Q(buf9[13]) );
  DFF_X1 \buf1_reg[12]  ( .D(element1[12]), .CK(clock), .Q(buf1[12]) );
  DFF_X1 \buf2_reg[12]  ( .D(buf1[12]), .CK(clock), .Q(buf2[12]) );
  DFF_X1 \buf3_reg[12]  ( .D(buf2[12]), .CK(clock), .Q(buf3[12]) );
  DFF_X1 \buf4_reg[12]  ( .D(buf3[12]), .CK(clock), .Q(buf4[12]) );
  DFF_X1 \buf5_reg[12]  ( .D(buf4[12]), .CK(clock), .Q(buf5[12]) );
  DFF_X1 \buf6_reg[12]  ( .D(buf5[12]), .CK(clock), .Q(buf6[12]) );
  DFF_X1 \buf7_reg[12]  ( .D(buf6[12]), .CK(clock), .Q(buf7[12]) );
  DFF_X1 \buf8_reg[12]  ( .D(buf7[12]), .CK(clock), .Q(buf8[12]) );
  DFF_X1 \buf9_reg[12]  ( .D(buf8[12]), .CK(clock), .Q(buf9[12]) );
  DFF_X1 \buf1_reg[11]  ( .D(element1[11]), .CK(clock), .Q(buf1[11]) );
  DFF_X1 \buf2_reg[11]  ( .D(buf1[11]), .CK(clock), .Q(buf2[11]) );
  DFF_X1 \buf3_reg[11]  ( .D(buf2[11]), .CK(clock), .Q(buf3[11]) );
  DFF_X1 \buf4_reg[11]  ( .D(buf3[11]), .CK(clock), .Q(buf4[11]) );
  DFF_X1 \buf5_reg[11]  ( .D(buf4[11]), .CK(clock), .Q(buf5[11]) );
  DFF_X1 \buf6_reg[11]  ( .D(buf5[11]), .CK(clock), .Q(buf6[11]) );
  DFF_X1 \buf7_reg[11]  ( .D(buf6[11]), .CK(clock), .Q(buf7[11]) );
  DFF_X1 \buf8_reg[11]  ( .D(buf7[11]), .CK(clock), .Q(buf8[11]) );
  DFF_X1 \buf9_reg[11]  ( .D(buf8[11]), .CK(clock), .Q(buf9[11]) );
  DFF_X1 \buf1_reg[10]  ( .D(element1[10]), .CK(clock), .Q(buf1[10]) );
  DFF_X1 \buf2_reg[10]  ( .D(buf1[10]), .CK(clock), .Q(buf2[10]) );
  DFF_X1 \buf3_reg[10]  ( .D(buf2[10]), .CK(clock), .Q(buf3[10]) );
  DFF_X1 \buf4_reg[10]  ( .D(buf3[10]), .CK(clock), .Q(buf4[10]) );
  DFF_X1 \buf5_reg[10]  ( .D(buf4[10]), .CK(clock), .Q(buf5[10]) );
  DFF_X1 \buf6_reg[10]  ( .D(buf5[10]), .CK(clock), .Q(buf6[10]) );
  DFF_X1 \buf7_reg[10]  ( .D(buf6[10]), .CK(clock), .Q(buf7[10]) );
  DFF_X1 \buf8_reg[10]  ( .D(buf7[10]), .CK(clock), .Q(buf8[10]) );
  DFF_X1 \buf9_reg[10]  ( .D(buf8[10]), .CK(clock), .Q(buf9[10]) );
  DFF_X1 \buf1_reg[9]  ( .D(element1[9]), .CK(clock), .Q(buf1[9]) );
  DFF_X1 \buf2_reg[9]  ( .D(buf1[9]), .CK(clock), .Q(buf2[9]) );
  DFF_X1 \buf3_reg[9]  ( .D(buf2[9]), .CK(clock), .Q(buf3[9]) );
  DFF_X1 \buf4_reg[9]  ( .D(buf3[9]), .CK(clock), .Q(buf4[9]) );
  DFF_X1 \buf5_reg[9]  ( .D(buf4[9]), .CK(clock), .Q(buf5[9]) );
  DFF_X1 \buf6_reg[9]  ( .D(buf5[9]), .CK(clock), .Q(buf6[9]) );
  DFF_X1 \buf7_reg[9]  ( .D(buf6[9]), .CK(clock), .Q(buf7[9]) );
  DFF_X1 \buf8_reg[9]  ( .D(buf7[9]), .CK(clock), .Q(buf8[9]) );
  DFF_X1 \buf9_reg[9]  ( .D(buf8[9]), .CK(clock), .Q(buf9[9]) );
  DFF_X1 \buf1_reg[8]  ( .D(element1[8]), .CK(clock), .Q(buf1[8]) );
  DFF_X1 \buf2_reg[8]  ( .D(buf1[8]), .CK(clock), .Q(buf2[8]) );
  DFF_X1 \buf3_reg[8]  ( .D(buf2[8]), .CK(clock), .Q(buf3[8]) );
  DFF_X1 \buf4_reg[8]  ( .D(buf3[8]), .CK(clock), .Q(buf4[8]) );
  DFF_X1 \buf5_reg[8]  ( .D(buf4[8]), .CK(clock), .Q(buf5[8]) );
  DFF_X1 \buf6_reg[8]  ( .D(buf5[8]), .CK(clock), .Q(buf6[8]) );
  DFF_X1 \buf7_reg[8]  ( .D(buf6[8]), .CK(clock), .Q(buf7[8]) );
  DFF_X1 \buf8_reg[8]  ( .D(buf7[8]), .CK(clock), .Q(buf8[8]) );
  DFF_X1 \buf9_reg[8]  ( .D(buf8[8]), .CK(clock), .Q(buf9[8]) );
  DFF_X1 \buf1_reg[7]  ( .D(element1[7]), .CK(clock), .Q(buf1[7]) );
  DFF_X1 \buf2_reg[7]  ( .D(buf1[7]), .CK(clock), .Q(buf2[7]) );
  DFF_X1 \buf3_reg[7]  ( .D(buf2[7]), .CK(clock), .Q(buf3[7]) );
  DFF_X1 \buf4_reg[7]  ( .D(buf3[7]), .CK(clock), .Q(buf4[7]) );
  DFF_X1 \buf5_reg[7]  ( .D(buf4[7]), .CK(clock), .Q(buf5[7]) );
  DFF_X1 \buf6_reg[7]  ( .D(buf5[7]), .CK(clock), .Q(buf6[7]) );
  DFF_X1 \buf7_reg[7]  ( .D(buf6[7]), .CK(clock), .Q(buf7[7]) );
  DFF_X1 \buf8_reg[7]  ( .D(buf7[7]), .CK(clock), .Q(buf8[7]) );
  DFF_X1 \buf9_reg[7]  ( .D(buf8[7]), .CK(clock), .Q(buf9[7]) );
  DFF_X1 \buf1_reg[6]  ( .D(element1[6]), .CK(clock), .Q(buf1[6]) );
  DFF_X1 \buf2_reg[6]  ( .D(buf1[6]), .CK(clock), .Q(buf2[6]) );
  DFF_X1 \buf3_reg[6]  ( .D(buf2[6]), .CK(clock), .Q(buf3[6]) );
  DFF_X1 \buf4_reg[6]  ( .D(buf3[6]), .CK(clock), .Q(buf4[6]) );
  DFF_X1 \buf5_reg[6]  ( .D(buf4[6]), .CK(clock), .Q(buf5[6]) );
  DFF_X1 \buf6_reg[6]  ( .D(buf5[6]), .CK(clock), .Q(buf6[6]) );
  DFF_X1 \buf7_reg[6]  ( .D(buf6[6]), .CK(clock), .Q(buf7[6]) );
  DFF_X1 \buf8_reg[6]  ( .D(buf7[6]), .CK(clock), .Q(buf8[6]) );
  DFF_X1 \buf9_reg[6]  ( .D(buf8[6]), .CK(clock), .Q(buf9[6]) );
  DFF_X1 \buf1_reg[5]  ( .D(element1[5]), .CK(clock), .Q(buf1[5]) );
  DFF_X1 \buf2_reg[5]  ( .D(buf1[5]), .CK(clock), .Q(buf2[5]) );
  DFF_X1 \buf3_reg[5]  ( .D(buf2[5]), .CK(clock), .Q(buf3[5]) );
  DFF_X1 \buf4_reg[5]  ( .D(buf3[5]), .CK(clock), .Q(buf4[5]) );
  DFF_X1 \buf5_reg[5]  ( .D(buf4[5]), .CK(clock), .Q(buf5[5]) );
  DFF_X1 \buf6_reg[5]  ( .D(buf5[5]), .CK(clock), .Q(buf6[5]) );
  DFF_X1 \buf7_reg[5]  ( .D(buf6[5]), .CK(clock), .Q(buf7[5]) );
  DFF_X1 \buf8_reg[5]  ( .D(buf7[5]), .CK(clock), .Q(buf8[5]) );
  DFF_X1 \buf9_reg[5]  ( .D(buf8[5]), .CK(clock), .Q(buf9[5]) );
  DFF_X1 \buf1_reg[4]  ( .D(element1[4]), .CK(clock), .Q(buf1[4]) );
  DFF_X1 \buf2_reg[4]  ( .D(buf1[4]), .CK(clock), .Q(buf2[4]) );
  DFF_X1 \buf3_reg[4]  ( .D(buf2[4]), .CK(clock), .Q(buf3[4]) );
  DFF_X1 \buf4_reg[4]  ( .D(buf3[4]), .CK(clock), .Q(buf4[4]) );
  DFF_X1 \buf5_reg[4]  ( .D(buf4[4]), .CK(clock), .Q(buf5[4]) );
  DFF_X1 \buf6_reg[4]  ( .D(buf5[4]), .CK(clock), .Q(buf6[4]) );
  DFF_X1 \buf7_reg[4]  ( .D(buf6[4]), .CK(clock), .Q(buf7[4]) );
  DFF_X1 \buf8_reg[4]  ( .D(buf7[4]), .CK(clock), .Q(buf8[4]) );
  DFF_X1 \buf9_reg[4]  ( .D(buf8[4]), .CK(clock), .Q(buf9[4]) );
  DFF_X1 \buf1_reg[3]  ( .D(element1[3]), .CK(clock), .Q(buf1[3]) );
  DFF_X1 \buf2_reg[3]  ( .D(buf1[3]), .CK(clock), .Q(buf2[3]) );
  DFF_X1 \buf3_reg[3]  ( .D(buf2[3]), .CK(clock), .Q(buf3[3]) );
  DFF_X1 \buf4_reg[3]  ( .D(buf3[3]), .CK(clock), .Q(buf4[3]) );
  DFF_X1 \buf5_reg[3]  ( .D(buf4[3]), .CK(clock), .Q(buf5[3]) );
  DFF_X1 \buf6_reg[3]  ( .D(buf5[3]), .CK(clock), .Q(buf6[3]) );
  DFF_X1 \buf7_reg[3]  ( .D(buf6[3]), .CK(clock), .Q(buf7[3]) );
  DFF_X1 \buf8_reg[3]  ( .D(buf7[3]), .CK(clock), .Q(buf8[3]) );
  DFF_X1 \buf9_reg[3]  ( .D(buf8[3]), .CK(clock), .Q(buf9[3]) );
  DFF_X1 \buf1_reg[2]  ( .D(element1[2]), .CK(clock), .Q(buf1[2]) );
  DFF_X1 \buf2_reg[2]  ( .D(buf1[2]), .CK(clock), .Q(buf2[2]) );
  DFF_X1 \buf3_reg[2]  ( .D(buf2[2]), .CK(clock), .Q(buf3[2]) );
  DFF_X1 \buf4_reg[2]  ( .D(buf3[2]), .CK(clock), .Q(buf4[2]) );
  DFF_X1 \buf5_reg[2]  ( .D(buf4[2]), .CK(clock), .Q(buf5[2]) );
  DFF_X1 \buf6_reg[2]  ( .D(buf5[2]), .CK(clock), .Q(buf6[2]) );
  DFF_X1 \buf7_reg[2]  ( .D(buf6[2]), .CK(clock), .Q(buf7[2]) );
  DFF_X1 \buf8_reg[2]  ( .D(buf7[2]), .CK(clock), .Q(buf8[2]) );
  DFF_X1 \buf9_reg[2]  ( .D(buf8[2]), .CK(clock), .Q(buf9[2]) );
  DFF_X1 \buf1_reg[1]  ( .D(element1[1]), .CK(clock), .Q(buf1[1]) );
  DFF_X1 \buf2_reg[1]  ( .D(buf1[1]), .CK(clock), .Q(buf2[1]) );
  DFF_X1 \buf3_reg[1]  ( .D(buf2[1]), .CK(clock), .Q(buf3[1]) );
  DFF_X1 \buf4_reg[1]  ( .D(buf3[1]), .CK(clock), .Q(buf4[1]) );
  DFF_X1 \buf5_reg[1]  ( .D(buf4[1]), .CK(clock), .Q(buf5[1]) );
  DFF_X1 \buf6_reg[1]  ( .D(buf5[1]), .CK(clock), .Q(buf6[1]) );
  DFF_X1 \buf7_reg[1]  ( .D(buf6[1]), .CK(clock), .Q(buf7[1]) );
  DFF_X1 \buf8_reg[1]  ( .D(buf7[1]), .CK(clock), .Q(buf8[1]) );
  DFF_X1 \buf9_reg[1]  ( .D(buf8[1]), .CK(clock), .Q(buf9[1]) );
  DFF_X1 \buf1_reg[0]  ( .D(element1[0]), .CK(clock), .Q(buf1[0]) );
  DFF_X1 \buf2_reg[0]  ( .D(buf1[0]), .CK(clock), .Q(buf2[0]) );
  DFF_X1 \buf3_reg[0]  ( .D(buf2[0]), .CK(clock), .Q(buf3[0]) );
  DFF_X1 \buf4_reg[0]  ( .D(buf3[0]), .CK(clock), .Q(buf4[0]) );
  DFF_X1 \buf5_reg[0]  ( .D(buf4[0]), .CK(clock), .Q(buf5[0]) );
  DFF_X1 \buf6_reg[0]  ( .D(buf5[0]), .CK(clock), .Q(buf6[0]) );
  DFF_X1 \buf7_reg[0]  ( .D(buf6[0]), .CK(clock), .Q(buf7[0]) );
  DFF_X1 \buf8_reg[0]  ( .D(buf7[0]), .CK(clock), .Q(buf8[0]) );
  DFF_X1 \buf9_reg[0]  ( .D(buf8[0]), .CK(clock), .Q(buf9[0]) );
  DFF_X2 \buf10_reg[0]  ( .D(buf9[0]), .CK(clock), .Q(op2[0]) );
  DFF_X2 \buf10_reg[1]  ( .D(buf9[1]), .CK(clock), .Q(op2[1]) );
  DFF_X2 \buf10_reg[2]  ( .D(buf9[2]), .CK(clock), .Q(op2[2]) );
  DFF_X2 \buf10_reg[3]  ( .D(buf9[3]), .CK(clock), .Q(op2[3]) );
  DFF_X2 \buf10_reg[4]  ( .D(buf9[4]), .CK(clock), .Q(op2[4]) );
  DFF_X2 \buf10_reg[5]  ( .D(buf9[5]), .CK(clock), .Q(op2[5]) );
  DFF_X2 \buf10_reg[6]  ( .D(buf9[6]), .CK(clock), .Q(op2[6]) );
  DFF_X2 \buf10_reg[7]  ( .D(buf9[7]), .CK(clock), .Q(op2[7]) );
  DFF_X2 \buf10_reg[8]  ( .D(buf9[8]), .CK(clock), .Q(op2[8]) );
  DFF_X2 \buf10_reg[9]  ( .D(buf9[9]), .CK(clock), .Q(op2[9]) );
  DFF_X2 \buf10_reg[10]  ( .D(buf9[10]), .CK(clock), .Q(op2[10]) );
  DFF_X2 \buf10_reg[11]  ( .D(buf9[11]), .CK(clock), .Q(op2[11]) );
  DFF_X2 \buf10_reg[12]  ( .D(buf9[12]), .CK(clock), .Q(op2[12]) );
  DFF_X2 \buf10_reg[13]  ( .D(buf9[13]), .CK(clock), .Q(op2[13]) );
  DFF_X2 \buf10_reg[14]  ( .D(buf9[14]), .CK(clock), .Q(op2[14]) );
  DFF_X2 \buf10_reg[15]  ( .D(buf9[15]), .CK(clock), .Q(op2[15]) );
  DFF_X2 \buf10_reg[16]  ( .D(buf9[16]), .CK(clock), .Q(op2[16]) );
  DFF_X2 \buf10_reg[17]  ( .D(buf9[17]), .CK(clock), .Q(op2[17]) );
  DFF_X2 \buf10_reg[18]  ( .D(buf9[18]), .CK(clock), .Q(op2[18]) );
  DFF_X2 \buf10_reg[19]  ( .D(buf9[19]), .CK(clock), .Q(op2[19]) );
  DFF_X2 \buf10_reg[20]  ( .D(buf9[20]), .CK(clock), .Q(op2[20]) );
  DFF_X2 \buf10_reg[21]  ( .D(buf9[21]), .CK(clock), .Q(op2[21]) );
  DFF_X2 \buf10_reg[22]  ( .D(buf9[22]), .CK(clock), .Q(op2[22]) );
  DFF_X2 \buf10_reg[23]  ( .D(buf9[23]), .CK(clock), .Q(op2[23]) );
  DFF_X2 \buf10_reg[24]  ( .D(buf9[24]), .CK(clock), .Q(op1[0]) );
  DFF_X2 \buf10_reg[25]  ( .D(buf9[25]), .CK(clock), .Q(op1[1]) );
  DFF_X2 \buf10_reg[26]  ( .D(buf9[26]), .CK(clock), .Q(op1[2]) );
  DFF_X2 \buf10_reg[27]  ( .D(buf9[27]), .CK(clock), .Q(op1[3]) );
  DFF_X2 \buf10_reg[28]  ( .D(buf9[28]), .CK(clock), .Q(op1[4]) );
  DFF_X2 \buf10_reg[29]  ( .D(buf9[29]), .CK(clock), .Q(op1[5]) );
  DFF_X2 \buf10_reg[30]  ( .D(buf9[30]), .CK(clock), .Q(op1[6]) );
  DFF_X2 \buf10_reg[31]  ( .D(buf9[31]), .CK(clock), .Q(op1[7]) );
  DFF_X2 \buf10_reg[32]  ( .D(buf9[32]), .CK(clock), .Q(op1[8]) );
  DFF_X2 \buf10_reg[33]  ( .D(buf9[33]), .CK(clock), .Q(op1[9]) );
  DFF_X2 \buf10_reg[34]  ( .D(buf9[34]), .CK(clock), .Q(op1[10]) );
  DFF_X2 \buf10_reg[35]  ( .D(buf9[35]), .CK(clock), .Q(op1[11]) );
  DFF_X2 \buf10_reg[36]  ( .D(buf9[36]), .CK(clock), .Q(op1[12]) );
  DFF_X2 \buf10_reg[37]  ( .D(buf9[37]), .CK(clock), .Q(op1[13]) );
  DFF_X2 \buf10_reg[38]  ( .D(buf9[38]), .CK(clock), .Q(op1[14]) );
  DFF_X2 \buf10_reg[39]  ( .D(buf9[39]), .CK(clock), .Q(op1[15]) );
  DFF_X2 \buf10_reg[40]  ( .D(buf9[40]), .CK(clock), .Q(op1[16]) );
  DFF_X2 \buf10_reg[41]  ( .D(buf9[41]), .CK(clock), .Q(op1[17]) );
  DFF_X2 \buf10_reg[42]  ( .D(buf9[42]), .CK(clock), .Q(op1[18]) );
  DFF_X2 \buf10_reg[43]  ( .D(buf9[43]), .CK(clock), .Q(op1[19]) );
  DFF_X2 \buf10_reg[44]  ( .D(buf9[44]), .CK(clock), .Q(op1[20]) );
  DFF_X2 \buf10_reg[45]  ( .D(buf9[45]), .CK(clock), .Q(op1[21]) );
  DFF_X2 \buf10_reg[46]  ( .D(buf9[46]), .CK(clock), .Q(op1[22]) );
  DFF_X2 \buf10_reg[47]  ( .D(buf9[47]), .CK(clock), .Q(op1[23]) );
endmodule


module syncMult ( clock, SyncY, SyncMultY, multinput, mult_output );
  input [48:0] SyncY;
  output [47:0] SyncMultY;
  input [47:0] multinput;
  output [48:0] mult_output;
  input clock;
  wire   bit_buf1, bit_buf2, bit_buf3, bit_buf4, bit_buf5, bit_buf6, bit_buf7,
         bit_buf8;

  DFF_X1 bit_buf1_reg ( .D(SyncY[48]), .CK(clock), .Q(bit_buf1) );
  DFF_X1 bit_buf2_reg ( .D(bit_buf1), .CK(clock), .Q(bit_buf2) );
  DFF_X1 bit_buf3_reg ( .D(bit_buf2), .CK(clock), .Q(bit_buf3) );
  DFF_X1 bit_buf4_reg ( .D(bit_buf3), .CK(clock), .Q(bit_buf4) );
  DFF_X1 bit_buf5_reg ( .D(bit_buf4), .CK(clock), .Q(bit_buf5) );
  DFF_X1 bit_buf6_reg ( .D(bit_buf5), .CK(clock), .Q(bit_buf6) );
  DFF_X1 bit_buf7_reg ( .D(bit_buf6), .CK(clock), .Q(bit_buf7) );
  DFF_X1 bit_buf8_reg ( .D(bit_buf7), .CK(clock), .Q(bit_buf8) );
  DFF_X2 bit_buf9_reg ( .D(bit_buf8), .CK(clock), .Q(mult_output[48]) );
  BUF_X4 U3 ( .A(multinput[6]), .Z(mult_output[6]) );
  BUF_X4 U4 ( .A(multinput[30]), .Z(mult_output[30]) );
  BUF_X4 U5 ( .A(multinput[31]), .Z(mult_output[31]) );
  BUF_X4 U6 ( .A(multinput[32]), .Z(mult_output[32]) );
  BUF_X4 U7 ( .A(multinput[9]), .Z(mult_output[9]) );
  BUF_X4 U8 ( .A(multinput[4]), .Z(mult_output[4]) );
  BUF_X4 U9 ( .A(multinput[10]), .Z(mult_output[10]) );
  BUF_X4 U10 ( .A(multinput[13]), .Z(mult_output[13]) );
  BUF_X4 U11 ( .A(multinput[16]), .Z(mult_output[16]) );
  BUF_X4 U12 ( .A(multinput[19]), .Z(mult_output[19]) );
  BUF_X4 U13 ( .A(multinput[21]), .Z(mult_output[21]) );
  BUF_X4 U14 ( .A(multinput[34]), .Z(mult_output[34]) );
  BUF_X4 U15 ( .A(multinput[37]), .Z(mult_output[37]) );
  BUF_X4 U16 ( .A(multinput[40]), .Z(mult_output[40]) );
  BUF_X4 U17 ( .A(multinput[43]), .Z(mult_output[43]) );
  BUF_X4 U18 ( .A(multinput[1]), .Z(mult_output[1]) );
  BUF_X4 U19 ( .A(multinput[2]), .Z(mult_output[2]) );
  BUF_X4 U20 ( .A(multinput[5]), .Z(mult_output[5]) );
  BUF_X4 U21 ( .A(multinput[11]), .Z(mult_output[11]) );
  BUF_X4 U22 ( .A(multinput[14]), .Z(mult_output[14]) );
  BUF_X4 U23 ( .A(multinput[17]), .Z(mult_output[17]) );
  BUF_X4 U24 ( .A(multinput[22]), .Z(mult_output[22]) );
  BUF_X4 U25 ( .A(multinput[0]), .Z(mult_output[0]) );
  BUF_X4 U26 ( .A(multinput[3]), .Z(mult_output[3]) );
  BUF_X4 U27 ( .A(multinput[7]), .Z(mult_output[7]) );
  BUF_X4 U28 ( .A(multinput[8]), .Z(mult_output[8]) );
  BUF_X4 U29 ( .A(multinput[12]), .Z(mult_output[12]) );
  BUF_X4 U30 ( .A(multinput[15]), .Z(mult_output[15]) );
  BUF_X4 U31 ( .A(multinput[18]), .Z(mult_output[18]) );
  BUF_X4 U32 ( .A(multinput[20]), .Z(mult_output[20]) );
  BUF_X4 U33 ( .A(multinput[23]), .Z(mult_output[23]) );
  BUF_X4 U34 ( .A(multinput[33]), .Z(mult_output[33]) );
  BUF_X4 U35 ( .A(multinput[28]), .Z(mult_output[28]) );
  BUF_X4 U36 ( .A(multinput[45]), .Z(mult_output[45]) );
  BUF_X4 U37 ( .A(multinput[24]), .Z(mult_output[24]) );
  BUF_X4 U38 ( .A(multinput[27]), .Z(mult_output[27]) );
  BUF_X4 U39 ( .A(multinput[36]), .Z(mult_output[36]) );
  BUF_X4 U40 ( .A(multinput[39]), .Z(mult_output[39]) );
  BUF_X4 U41 ( .A(multinput[42]), .Z(mult_output[42]) );
  BUF_X4 U42 ( .A(multinput[44]), .Z(mult_output[44]) );
  BUF_X4 U43 ( .A(multinput[47]), .Z(mult_output[47]) );
  BUF_X4 U44 ( .A(multinput[25]), .Z(mult_output[25]) );
  BUF_X4 U45 ( .A(multinput[26]), .Z(mult_output[26]) );
  BUF_X4 U46 ( .A(multinput[29]), .Z(mult_output[29]) );
  BUF_X4 U47 ( .A(multinput[35]), .Z(mult_output[35]) );
  BUF_X4 U48 ( .A(multinput[38]), .Z(mult_output[38]) );
  BUF_X4 U49 ( .A(multinput[41]), .Z(mult_output[41]) );
  BUF_X4 U50 ( .A(multinput[46]), .Z(mult_output[46]) );
  BUF_X4 U51 ( .A(SyncY[0]), .Z(SyncMultY[0]) );
  BUF_X4 U52 ( .A(SyncY[1]), .Z(SyncMultY[1]) );
  BUF_X4 U53 ( .A(SyncY[2]), .Z(SyncMultY[2]) );
  BUF_X4 U54 ( .A(SyncY[3]), .Z(SyncMultY[3]) );
  BUF_X4 U55 ( .A(SyncY[4]), .Z(SyncMultY[4]) );
  BUF_X4 U56 ( .A(SyncY[5]), .Z(SyncMultY[5]) );
  BUF_X4 U57 ( .A(SyncY[6]), .Z(SyncMultY[6]) );
  BUF_X4 U58 ( .A(SyncY[7]), .Z(SyncMultY[7]) );
  BUF_X4 U59 ( .A(SyncY[8]), .Z(SyncMultY[8]) );
  BUF_X4 U60 ( .A(SyncY[9]), .Z(SyncMultY[9]) );
  BUF_X4 U61 ( .A(SyncY[10]), .Z(SyncMultY[10]) );
  BUF_X4 U62 ( .A(SyncY[11]), .Z(SyncMultY[11]) );
  BUF_X4 U63 ( .A(SyncY[12]), .Z(SyncMultY[12]) );
  BUF_X4 U64 ( .A(SyncY[13]), .Z(SyncMultY[13]) );
  BUF_X4 U65 ( .A(SyncY[14]), .Z(SyncMultY[14]) );
  BUF_X4 U66 ( .A(SyncY[15]), .Z(SyncMultY[15]) );
  BUF_X4 U67 ( .A(SyncY[16]), .Z(SyncMultY[16]) );
  BUF_X4 U68 ( .A(SyncY[17]), .Z(SyncMultY[17]) );
  BUF_X4 U69 ( .A(SyncY[18]), .Z(SyncMultY[18]) );
  BUF_X4 U70 ( .A(SyncY[19]), .Z(SyncMultY[19]) );
  BUF_X4 U71 ( .A(SyncY[20]), .Z(SyncMultY[20]) );
  BUF_X4 U72 ( .A(SyncY[21]), .Z(SyncMultY[21]) );
  BUF_X4 U73 ( .A(SyncY[22]), .Z(SyncMultY[22]) );
  BUF_X4 U74 ( .A(SyncY[23]), .Z(SyncMultY[23]) );
  BUF_X4 U75 ( .A(SyncY[24]), .Z(SyncMultY[24]) );
  BUF_X4 U76 ( .A(SyncY[25]), .Z(SyncMultY[25]) );
  BUF_X4 U77 ( .A(SyncY[26]), .Z(SyncMultY[26]) );
  BUF_X4 U78 ( .A(SyncY[27]), .Z(SyncMultY[27]) );
  BUF_X4 U79 ( .A(SyncY[28]), .Z(SyncMultY[28]) );
  BUF_X4 U80 ( .A(SyncY[29]), .Z(SyncMultY[29]) );
  BUF_X4 U81 ( .A(SyncY[30]), .Z(SyncMultY[30]) );
  BUF_X4 U82 ( .A(SyncY[31]), .Z(SyncMultY[31]) );
  BUF_X4 U83 ( .A(SyncY[32]), .Z(SyncMultY[32]) );
  BUF_X4 U84 ( .A(SyncY[33]), .Z(SyncMultY[33]) );
  BUF_X4 U85 ( .A(SyncY[34]), .Z(SyncMultY[34]) );
  BUF_X4 U86 ( .A(SyncY[35]), .Z(SyncMultY[35]) );
  BUF_X4 U87 ( .A(SyncY[36]), .Z(SyncMultY[36]) );
  BUF_X4 U88 ( .A(SyncY[37]), .Z(SyncMultY[37]) );
  BUF_X4 U89 ( .A(SyncY[38]), .Z(SyncMultY[38]) );
  BUF_X4 U90 ( .A(SyncY[39]), .Z(SyncMultY[39]) );
  BUF_X4 U91 ( .A(SyncY[40]), .Z(SyncMultY[40]) );
  BUF_X4 U92 ( .A(SyncY[41]), .Z(SyncMultY[41]) );
  BUF_X4 U93 ( .A(SyncY[42]), .Z(SyncMultY[42]) );
  BUF_X4 U94 ( .A(SyncY[43]), .Z(SyncMultY[43]) );
  BUF_X4 U95 ( .A(SyncY[44]), .Z(SyncMultY[44]) );
  BUF_X4 U96 ( .A(SyncY[45]), .Z(SyncMultY[45]) );
  BUF_X4 U97 ( .A(SyncY[47]), .Z(SyncMultY[47]) );
  BUF_X4 U98 ( .A(SyncY[46]), .Z(SyncMultY[46]) );
endmodule


module controller2_1 ( clock, reset, accum_in, feedback, set_bit, count, 
        count2, element, adder_out1, adder_out2, adder_out3, adder_out4 );
  input [24:0] accum_in;
  output [23:0] feedback;
  output [4:0] count;
  output [2:0] count2;
  input [24:0] element;
  output [23:0] adder_out1;
  output [23:0] adder_out2;
  output [23:0] adder_out3;
  output [23:0] adder_out4;
  input clock, reset, set_bit;
  wire   N7, N8, N9, N10, N11, N12, N13, N14, N24, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, \add_32/carry[4] ,
         \add_32/carry[3] , \add_32/carry[2] , n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576;

  DFF_X1 \count_reg[0]  ( .D(N11), .CK(clock), .Q(count[0]), .QN(n549) );
  DFF_X1 \count_reg[1]  ( .D(N12), .CK(clock), .Q(count[1]), .QN(n548) );
  DFF_X1 \count_reg[2]  ( .D(N13), .CK(clock), .Q(count[2]) );
  DFF_X1 \count_reg[3]  ( .D(N14), .CK(clock), .Q(count[3]) );
  DFF_X1 \count_reg[4]  ( .D(n44), .CK(clock), .Q(count[4]) );
  NOR2_X2 U101 ( .A1(n31), .A2(n567), .ZN(feedback[9]) );
  NOR2_X2 U102 ( .A1(n31), .A2(n568), .ZN(feedback[8]) );
  NOR2_X2 U103 ( .A1(n31), .A2(n569), .ZN(feedback[7]) );
  NOR2_X2 U104 ( .A1(n31), .A2(n570), .ZN(feedback[6]) );
  NOR2_X2 U105 ( .A1(n31), .A2(n571), .ZN(feedback[5]) );
  NOR2_X2 U106 ( .A1(n31), .A2(n572), .ZN(feedback[4]) );
  NOR2_X2 U107 ( .A1(n31), .A2(n573), .ZN(feedback[3]) );
  NOR2_X2 U108 ( .A1(n31), .A2(n574), .ZN(feedback[2]) );
  NOR2_X2 U109 ( .A1(n31), .A2(n553), .ZN(feedback[23]) );
  NOR2_X2 U110 ( .A1(n31), .A2(n554), .ZN(feedback[22]) );
  NOR2_X2 U111 ( .A1(n31), .A2(n555), .ZN(feedback[21]) );
  NOR2_X2 U112 ( .A1(n31), .A2(n556), .ZN(feedback[20]) );
  NOR2_X2 U113 ( .A1(n31), .A2(n575), .ZN(feedback[1]) );
  NOR2_X2 U114 ( .A1(n31), .A2(n557), .ZN(feedback[19]) );
  NOR2_X2 U115 ( .A1(n31), .A2(n558), .ZN(feedback[18]) );
  NOR2_X2 U116 ( .A1(n31), .A2(n559), .ZN(feedback[17]) );
  NOR2_X2 U117 ( .A1(n31), .A2(n560), .ZN(feedback[16]) );
  NOR2_X2 U118 ( .A1(n31), .A2(n561), .ZN(feedback[15]) );
  NOR2_X2 U119 ( .A1(n31), .A2(n562), .ZN(feedback[14]) );
  NOR2_X2 U120 ( .A1(n31), .A2(n563), .ZN(feedback[13]) );
  NOR2_X2 U121 ( .A1(n31), .A2(n564), .ZN(feedback[12]) );
  NOR2_X2 U122 ( .A1(n31), .A2(n565), .ZN(feedback[11]) );
  NOR2_X2 U123 ( .A1(n31), .A2(n566), .ZN(feedback[10]) );
  NOR2_X2 U124 ( .A1(n31), .A2(n576), .ZN(feedback[0]) );
  NAND2_X2 U125 ( .A1(N24), .A2(n552), .ZN(n31) );
  NOR2_X2 U127 ( .A1(set_bit), .A2(reset), .ZN(n35) );
  NAND4_X2 U128 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n34) );
  NOR3_X2 U129 ( .A1(element[18]), .A2(element[1]), .A3(element[19]), .ZN(n39)
         );
  NOR3_X2 U130 ( .A1(element[15]), .A2(element[17]), .A3(element[16]), .ZN(n38) );
  NOR3_X2 U131 ( .A1(element[12]), .A2(element[14]), .A3(element[13]), .ZN(n37) );
  NOR3_X2 U132 ( .A1(element[0]), .A2(element[11]), .A3(element[10]), .ZN(n36)
         );
  NAND4_X2 U133 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n33) );
  NOR4_X2 U134 ( .A1(element[9]), .A2(element[8]), .A3(element[7]), .A4(
        element[6]), .ZN(n43) );
  NOR3_X2 U135 ( .A1(element[3]), .A2(element[5]), .A3(element[4]), .ZN(n42)
         );
  NOR3_X2 U136 ( .A1(element[23]), .A2(element[2]), .A3(element[24]), .ZN(n41)
         );
  NOR3_X2 U137 ( .A1(element[20]), .A2(element[22]), .A3(element[21]), .ZN(n40) );
  AND2_X1 U164 ( .A1(N10), .A2(n551), .ZN(n44) );
  AND2_X1 U165 ( .A1(N9), .A2(n551), .ZN(N14) );
  AND2_X1 U166 ( .A1(N8), .A2(n551), .ZN(N13) );
  AND2_X1 U167 ( .A1(N7), .A2(n551), .ZN(N12) );
  HA_X1 \add_32/U1_1_1  ( .A(count[1]), .B(count[0]), .CO(\add_32/carry[2] ), 
        .S(N7) );
  HA_X1 \add_32/U1_1_2  ( .A(count[2]), .B(\add_32/carry[2] ), .CO(
        \add_32/carry[3] ), .S(N8) );
  HA_X1 \add_32/U1_1_3  ( .A(count[3]), .B(\add_32/carry[3] ), .CO(
        \add_32/carry[4] ), .S(N9) );
  INV_X4 U5 ( .A(1'b1), .ZN(adder_out4[0]) );
  INV_X4 U126 ( .A(1'b1), .ZN(adder_out4[1]) );
  INV_X4 U139 ( .A(1'b1), .ZN(adder_out4[2]) );
  INV_X4 U141 ( .A(1'b1), .ZN(adder_out4[3]) );
  INV_X4 U143 ( .A(1'b1), .ZN(adder_out4[4]) );
  INV_X4 U145 ( .A(1'b1), .ZN(adder_out4[5]) );
  INV_X4 U147 ( .A(1'b1), .ZN(adder_out4[6]) );
  INV_X4 U149 ( .A(1'b1), .ZN(adder_out4[7]) );
  INV_X4 U151 ( .A(1'b1), .ZN(adder_out4[8]) );
  INV_X4 U153 ( .A(1'b1), .ZN(adder_out4[9]) );
  INV_X4 U155 ( .A(1'b1), .ZN(adder_out4[10]) );
  INV_X4 U157 ( .A(1'b1), .ZN(adder_out4[11]) );
  INV_X4 U159 ( .A(1'b1), .ZN(adder_out4[12]) );
  INV_X4 U161 ( .A(1'b1), .ZN(adder_out4[13]) );
  INV_X4 U163 ( .A(1'b1), .ZN(adder_out4[14]) );
  INV_X4 U169 ( .A(1'b1), .ZN(adder_out4[15]) );
  INV_X4 U171 ( .A(1'b1), .ZN(adder_out4[16]) );
  INV_X4 U173 ( .A(1'b1), .ZN(adder_out4[17]) );
  INV_X4 U175 ( .A(1'b1), .ZN(adder_out4[18]) );
  INV_X4 U177 ( .A(1'b1), .ZN(adder_out4[19]) );
  INV_X4 U179 ( .A(1'b1), .ZN(adder_out4[20]) );
  INV_X4 U181 ( .A(1'b1), .ZN(adder_out4[21]) );
  INV_X4 U183 ( .A(1'b1), .ZN(adder_out4[22]) );
  INV_X4 U185 ( .A(1'b1), .ZN(adder_out4[23]) );
  INV_X4 U187 ( .A(1'b1), .ZN(adder_out3[0]) );
  INV_X4 U189 ( .A(1'b1), .ZN(adder_out3[1]) );
  INV_X4 U191 ( .A(1'b1), .ZN(adder_out3[2]) );
  INV_X4 U193 ( .A(1'b1), .ZN(adder_out3[3]) );
  INV_X4 U195 ( .A(1'b1), .ZN(adder_out3[4]) );
  INV_X4 U197 ( .A(1'b1), .ZN(adder_out3[5]) );
  INV_X4 U199 ( .A(1'b1), .ZN(adder_out3[6]) );
  INV_X4 U201 ( .A(1'b1), .ZN(adder_out3[7]) );
  INV_X4 U203 ( .A(1'b1), .ZN(adder_out3[8]) );
  INV_X4 U205 ( .A(1'b1), .ZN(adder_out3[9]) );
  INV_X4 U207 ( .A(1'b1), .ZN(adder_out3[10]) );
  INV_X4 U209 ( .A(1'b1), .ZN(adder_out3[11]) );
  INV_X4 U211 ( .A(1'b1), .ZN(adder_out3[12]) );
  INV_X4 U213 ( .A(1'b1), .ZN(adder_out3[13]) );
  INV_X4 U215 ( .A(1'b1), .ZN(adder_out3[14]) );
  INV_X4 U217 ( .A(1'b1), .ZN(adder_out3[15]) );
  INV_X4 U219 ( .A(1'b1), .ZN(adder_out3[16]) );
  INV_X4 U221 ( .A(1'b1), .ZN(adder_out3[17]) );
  INV_X4 U223 ( .A(1'b1), .ZN(adder_out3[18]) );
  INV_X4 U225 ( .A(1'b1), .ZN(adder_out3[19]) );
  INV_X4 U227 ( .A(1'b1), .ZN(adder_out3[20]) );
  INV_X4 U229 ( .A(1'b1), .ZN(adder_out3[21]) );
  INV_X4 U231 ( .A(1'b1), .ZN(adder_out3[22]) );
  INV_X4 U233 ( .A(1'b1), .ZN(adder_out3[23]) );
  INV_X4 U235 ( .A(1'b1), .ZN(adder_out2[0]) );
  INV_X4 U237 ( .A(1'b1), .ZN(adder_out2[1]) );
  INV_X4 U239 ( .A(1'b1), .ZN(adder_out2[2]) );
  INV_X4 U241 ( .A(1'b1), .ZN(adder_out2[3]) );
  INV_X4 U243 ( .A(1'b1), .ZN(adder_out2[4]) );
  INV_X4 U245 ( .A(1'b1), .ZN(adder_out2[5]) );
  INV_X4 U247 ( .A(1'b1), .ZN(adder_out2[6]) );
  INV_X4 U249 ( .A(1'b1), .ZN(adder_out2[7]) );
  INV_X4 U251 ( .A(1'b1), .ZN(adder_out2[8]) );
  INV_X4 U253 ( .A(1'b1), .ZN(adder_out2[9]) );
  INV_X4 U255 ( .A(1'b1), .ZN(adder_out2[10]) );
  INV_X4 U257 ( .A(1'b1), .ZN(adder_out2[11]) );
  INV_X4 U259 ( .A(1'b1), .ZN(adder_out2[12]) );
  INV_X4 U261 ( .A(1'b1), .ZN(adder_out2[13]) );
  INV_X4 U263 ( .A(1'b1), .ZN(adder_out2[14]) );
  INV_X4 U265 ( .A(1'b1), .ZN(adder_out2[15]) );
  INV_X4 U267 ( .A(1'b1), .ZN(adder_out2[16]) );
  INV_X4 U269 ( .A(1'b1), .ZN(adder_out2[17]) );
  INV_X4 U271 ( .A(1'b1), .ZN(adder_out2[18]) );
  INV_X4 U273 ( .A(1'b1), .ZN(adder_out2[19]) );
  INV_X4 U275 ( .A(1'b1), .ZN(adder_out2[20]) );
  INV_X4 U277 ( .A(1'b1), .ZN(adder_out2[21]) );
  INV_X4 U279 ( .A(1'b1), .ZN(adder_out2[22]) );
  INV_X4 U281 ( .A(1'b1), .ZN(adder_out2[23]) );
  INV_X4 U283 ( .A(1'b1), .ZN(adder_out1[0]) );
  INV_X4 U285 ( .A(1'b1), .ZN(adder_out1[1]) );
  INV_X4 U287 ( .A(1'b1), .ZN(adder_out1[2]) );
  INV_X4 U289 ( .A(1'b1), .ZN(adder_out1[3]) );
  INV_X4 U291 ( .A(1'b1), .ZN(adder_out1[4]) );
  INV_X4 U293 ( .A(1'b1), .ZN(adder_out1[5]) );
  INV_X4 U295 ( .A(1'b1), .ZN(adder_out1[6]) );
  INV_X4 U297 ( .A(1'b1), .ZN(adder_out1[7]) );
  INV_X4 U299 ( .A(1'b1), .ZN(adder_out1[8]) );
  INV_X4 U301 ( .A(1'b1), .ZN(adder_out1[9]) );
  INV_X4 U303 ( .A(1'b1), .ZN(adder_out1[10]) );
  INV_X4 U305 ( .A(1'b1), .ZN(adder_out1[11]) );
  INV_X4 U307 ( .A(1'b1), .ZN(adder_out1[12]) );
  INV_X4 U309 ( .A(1'b1), .ZN(adder_out1[13]) );
  INV_X4 U311 ( .A(1'b1), .ZN(adder_out1[14]) );
  INV_X4 U313 ( .A(1'b1), .ZN(adder_out1[15]) );
  INV_X4 U315 ( .A(1'b1), .ZN(adder_out1[16]) );
  INV_X4 U317 ( .A(1'b1), .ZN(adder_out1[17]) );
  INV_X4 U319 ( .A(1'b1), .ZN(adder_out1[18]) );
  INV_X4 U321 ( .A(1'b1), .ZN(adder_out1[19]) );
  INV_X4 U323 ( .A(1'b1), .ZN(adder_out1[20]) );
  INV_X4 U325 ( .A(1'b1), .ZN(adder_out1[21]) );
  INV_X4 U327 ( .A(1'b1), .ZN(adder_out1[22]) );
  INV_X4 U329 ( .A(1'b1), .ZN(adder_out1[23]) );
  NOR2_X2 U331 ( .A1(n548), .A2(n549), .ZN(n550) );
  NOR2_X2 U332 ( .A1(count[0]), .A2(n32), .ZN(N11) );
  OAI21_X2 U333 ( .B1(n33), .B2(n34), .A(n35), .ZN(n32) );
  XOR2_X1 U334 ( .A(\add_32/carry[4] ), .B(count[4]), .Z(N10) );
  OR4_X1 U335 ( .A1(count[2]), .A2(n550), .A3(count[4]), .A4(count[3]), .ZN(
        N24) );
  INV_X4 U336 ( .A(n32), .ZN(n551) );
  INV_X4 U337 ( .A(set_bit), .ZN(n552) );
  INV_X4 U338 ( .A(accum_in[23]), .ZN(n553) );
  INV_X4 U339 ( .A(accum_in[22]), .ZN(n554) );
  INV_X4 U340 ( .A(accum_in[21]), .ZN(n555) );
  INV_X4 U341 ( .A(accum_in[20]), .ZN(n556) );
  INV_X4 U342 ( .A(accum_in[19]), .ZN(n557) );
  INV_X4 U343 ( .A(accum_in[18]), .ZN(n558) );
  INV_X4 U344 ( .A(accum_in[17]), .ZN(n559) );
  INV_X4 U345 ( .A(accum_in[16]), .ZN(n560) );
  INV_X4 U346 ( .A(accum_in[15]), .ZN(n561) );
  INV_X4 U347 ( .A(accum_in[14]), .ZN(n562) );
  INV_X4 U348 ( .A(accum_in[13]), .ZN(n563) );
  INV_X4 U349 ( .A(accum_in[12]), .ZN(n564) );
  INV_X4 U350 ( .A(accum_in[11]), .ZN(n565) );
  INV_X4 U351 ( .A(accum_in[10]), .ZN(n566) );
  INV_X4 U352 ( .A(accum_in[9]), .ZN(n567) );
  INV_X4 U353 ( .A(accum_in[8]), .ZN(n568) );
  INV_X4 U354 ( .A(accum_in[7]), .ZN(n569) );
  INV_X4 U355 ( .A(accum_in[6]), .ZN(n570) );
  INV_X4 U356 ( .A(accum_in[5]), .ZN(n571) );
  INV_X4 U357 ( .A(accum_in[4]), .ZN(n572) );
  INV_X4 U358 ( .A(accum_in[3]), .ZN(n573) );
  INV_X4 U359 ( .A(accum_in[2]), .ZN(n574) );
  INV_X4 U360 ( .A(accum_in[1]), .ZN(n575) );
  INV_X4 U361 ( .A(accum_in[0]), .ZN(n576) );
endmodule


module syncAccum_0 ( clock, mult_output, accum_input, accum_output, 
        accum_output25 );
  input [24:0] mult_output;
  output [23:0] accum_input;
  input [23:0] accum_output;
  output [24:0] accum_output25;
  input clock;
  wire   dirtybuff1, dirtybuff2, dirtybuff3;

  DFF_X1 dirtybuff1_reg ( .D(mult_output[24]), .CK(clock), .Q(dirtybuff1) );
  DFF_X1 dirtybuff2_reg ( .D(dirtybuff1), .CK(clock), .Q(dirtybuff2) );
  DFF_X1 dirtybuff3_reg ( .D(dirtybuff2), .CK(clock), .Q(dirtybuff3) );
  DFF_X1 dirtybuff4_reg ( .D(dirtybuff3), .CK(clock), .Q(accum_output25[24])
         );
  BUF_X4 U3 ( .A(mult_output[0]), .Z(accum_input[0]) );
  BUF_X4 U4 ( .A(mult_output[1]), .Z(accum_input[1]) );
  BUF_X4 U5 ( .A(mult_output[2]), .Z(accum_input[2]) );
  BUF_X4 U6 ( .A(mult_output[3]), .Z(accum_input[3]) );
  BUF_X4 U7 ( .A(mult_output[4]), .Z(accum_input[4]) );
  BUF_X4 U8 ( .A(mult_output[5]), .Z(accum_input[5]) );
  BUF_X4 U9 ( .A(mult_output[6]), .Z(accum_input[6]) );
  BUF_X4 U10 ( .A(mult_output[7]), .Z(accum_input[7]) );
  BUF_X4 U11 ( .A(mult_output[8]), .Z(accum_input[8]) );
  BUF_X4 U12 ( .A(mult_output[9]), .Z(accum_input[9]) );
  BUF_X4 U13 ( .A(mult_output[10]), .Z(accum_input[10]) );
  BUF_X4 U14 ( .A(mult_output[11]), .Z(accum_input[11]) );
  BUF_X4 U15 ( .A(mult_output[12]), .Z(accum_input[12]) );
  BUF_X4 U16 ( .A(mult_output[13]), .Z(accum_input[13]) );
  BUF_X4 U17 ( .A(mult_output[14]), .Z(accum_input[14]) );
  BUF_X4 U18 ( .A(mult_output[15]), .Z(accum_input[15]) );
  BUF_X4 U19 ( .A(mult_output[16]), .Z(accum_input[16]) );
  BUF_X4 U20 ( .A(mult_output[17]), .Z(accum_input[17]) );
  BUF_X4 U21 ( .A(mult_output[18]), .Z(accum_input[18]) );
  BUF_X4 U22 ( .A(mult_output[19]), .Z(accum_input[19]) );
  BUF_X4 U23 ( .A(mult_output[20]), .Z(accum_input[20]) );
  BUF_X4 U24 ( .A(mult_output[21]), .Z(accum_input[21]) );
  BUF_X4 U25 ( .A(mult_output[22]), .Z(accum_input[22]) );
  BUF_X4 U26 ( .A(mult_output[23]), .Z(accum_input[23]) );
  BUF_X4 U27 ( .A(accum_output[0]), .Z(accum_output25[0]) );
  BUF_X4 U28 ( .A(accum_output[1]), .Z(accum_output25[1]) );
  BUF_X4 U29 ( .A(accum_output[2]), .Z(accum_output25[2]) );
  BUF_X4 U30 ( .A(accum_output[3]), .Z(accum_output25[3]) );
  BUF_X4 U31 ( .A(accum_output[4]), .Z(accum_output25[4]) );
  BUF_X4 U32 ( .A(accum_output[5]), .Z(accum_output25[5]) );
  BUF_X4 U33 ( .A(accum_output[6]), .Z(accum_output25[6]) );
  BUF_X4 U34 ( .A(accum_output[7]), .Z(accum_output25[7]) );
  BUF_X4 U35 ( .A(accum_output[8]), .Z(accum_output25[8]) );
  BUF_X4 U36 ( .A(accum_output[9]), .Z(accum_output25[9]) );
  BUF_X4 U37 ( .A(accum_output[10]), .Z(accum_output25[10]) );
  BUF_X4 U38 ( .A(accum_output[11]), .Z(accum_output25[11]) );
  BUF_X4 U39 ( .A(accum_output[12]), .Z(accum_output25[12]) );
  BUF_X4 U40 ( .A(accum_output[13]), .Z(accum_output25[13]) );
  BUF_X4 U41 ( .A(accum_output[14]), .Z(accum_output25[14]) );
  BUF_X4 U42 ( .A(accum_output[15]), .Z(accum_output25[15]) );
  BUF_X4 U43 ( .A(accum_output[16]), .Z(accum_output25[16]) );
  BUF_X4 U44 ( .A(accum_output[17]), .Z(accum_output25[17]) );
  BUF_X4 U45 ( .A(accum_output[18]), .Z(accum_output25[18]) );
  BUF_X4 U46 ( .A(accum_output[19]), .Z(accum_output25[19]) );
  BUF_X4 U47 ( .A(accum_output[20]), .Z(accum_output25[20]) );
  BUF_X4 U48 ( .A(accum_output[21]), .Z(accum_output25[21]) );
  BUF_X4 U49 ( .A(accum_output[22]), .Z(accum_output25[22]) );
  BUF_X4 U50 ( .A(accum_output[23]), .Z(accum_output25[23]) );
endmodule


module controller2_0 ( clock, reset, accum_in, feedback, set_bit, count, 
        count2, element, adder_out1, adder_out2, adder_out3, adder_out4 );
  input [24:0] accum_in;
  output [23:0] feedback;
  output [4:0] count;
  output [2:0] count2;
  input [24:0] element;
  output [23:0] adder_out1;
  output [23:0] adder_out2;
  output [23:0] adder_out3;
  output [23:0] adder_out4;
  input clock, reset, set_bit;
  wire   \U10/Z_0 , \U10/Z_1 , \U10/Z_2 , \U10/Z_3 , \U10/Z_4 , \U10/Z_5 ,
         \U10/Z_6 , \U10/Z_7 , \U10/Z_8 , \U10/Z_9 , \U10/Z_10 , \U10/Z_11 ,
         \U10/Z_12 , \U10/Z_13 , \U10/Z_14 , \U10/Z_15 , \U10/Z_16 ,
         \U10/Z_17 , \U10/Z_18 , \U10/Z_19 , \U10/Z_20 , \U10/Z_21 ,
         \U10/Z_22 , \U10/Z_23 , \U10/DATA2_0 , \U10/DATA2_1 , \U10/DATA2_2 ,
         \U10/DATA2_3 , \U10/DATA2_4 , \U10/DATA2_5 , \U10/DATA2_6 ,
         \U10/DATA2_7 , \U10/DATA2_8 , \U10/DATA2_9 , \U10/DATA2_10 ,
         \U10/DATA2_11 , \U10/DATA2_12 , \U10/DATA2_13 , \U10/DATA2_14 ,
         \U10/DATA2_15 , \U10/DATA2_16 , \U10/DATA2_17 , \U10/DATA2_18 ,
         \U10/DATA2_19 , \U10/DATA2_20 , \U10/DATA2_21 , \U10/DATA2_22 ,
         \U10/DATA2_23 , \U4/Z_0 , \U4/Z_1 , \U4/Z_2 , \U4/Z_3 , \U4/DATA2_1 ,
         \U4/DATA2_2 , \U4/DATA2_3 , \add_32/carry[4] , \add_32/carry[3] ,
         \add_32/carry[2] , \add_32/A[0] , \add_32/A[1] , \add_32/A[2] ,
         \add_32/A[3] , \add_32/A[4] , n1, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576;
  assign feedback[0] = \U10/Z_0 ;
  assign feedback[1] = \U10/Z_1 ;
  assign feedback[2] = \U10/Z_2 ;
  assign feedback[3] = \U10/Z_3 ;
  assign feedback[4] = \U10/Z_4 ;
  assign feedback[5] = \U10/Z_5 ;
  assign feedback[6] = \U10/Z_6 ;
  assign feedback[7] = \U10/Z_7 ;
  assign feedback[8] = \U10/Z_8 ;
  assign feedback[9] = \U10/Z_9 ;
  assign feedback[10] = \U10/Z_10 ;
  assign feedback[11] = \U10/Z_11 ;
  assign feedback[12] = \U10/Z_12 ;
  assign feedback[13] = \U10/Z_13 ;
  assign feedback[14] = \U10/Z_14 ;
  assign feedback[15] = \U10/Z_15 ;
  assign feedback[16] = \U10/Z_16 ;
  assign feedback[17] = \U10/Z_17 ;
  assign feedback[18] = \U10/Z_18 ;
  assign feedback[19] = \U10/Z_19 ;
  assign feedback[20] = \U10/Z_20 ;
  assign feedback[21] = \U10/Z_21 ;
  assign feedback[22] = \U10/Z_22 ;
  assign feedback[23] = \U10/Z_23 ;
  assign \U10/DATA2_0  = accum_in[0];
  assign \U10/DATA2_1  = accum_in[1];
  assign \U10/DATA2_2  = accum_in[2];
  assign \U10/DATA2_3  = accum_in[3];
  assign \U10/DATA2_4  = accum_in[4];
  assign \U10/DATA2_5  = accum_in[5];
  assign \U10/DATA2_6  = accum_in[6];
  assign \U10/DATA2_7  = accum_in[7];
  assign \U10/DATA2_8  = accum_in[8];
  assign \U10/DATA2_9  = accum_in[9];
  assign \U10/DATA2_10  = accum_in[10];
  assign \U10/DATA2_11  = accum_in[11];
  assign \U10/DATA2_12  = accum_in[12];
  assign \U10/DATA2_13  = accum_in[13];
  assign \U10/DATA2_14  = accum_in[14];
  assign \U10/DATA2_15  = accum_in[15];
  assign \U10/DATA2_16  = accum_in[16];
  assign \U10/DATA2_17  = accum_in[17];
  assign \U10/DATA2_18  = accum_in[18];
  assign \U10/DATA2_19  = accum_in[19];
  assign \U10/DATA2_20  = accum_in[20];
  assign \U10/DATA2_21  = accum_in[21];
  assign \U10/DATA2_22  = accum_in[22];
  assign \U10/DATA2_23  = accum_in[23];
  assign count[0] = \add_32/A[0] ;
  assign count[1] = \add_32/A[1] ;
  assign count[2] = \add_32/A[2] ;
  assign count[3] = \add_32/A[3] ;
  assign count[4] = \add_32/A[4] ;

  HA_X1 \add_32/U1_1_1  ( .A(\add_32/A[1] ), .B(\add_32/A[0] ), .CO(
        \add_32/carry[2] ), .S(\U4/DATA2_1 ) );
  HA_X1 \add_32/U1_1_2  ( .A(\add_32/A[2] ), .B(\add_32/carry[2] ), .CO(
        \add_32/carry[3] ), .S(\U4/DATA2_2 ) );
  HA_X1 \add_32/U1_1_3  ( .A(\add_32/A[3] ), .B(\add_32/carry[3] ), .CO(
        \add_32/carry[4] ), .S(\U4/DATA2_3 ) );
  DFF_X1 \count_reg[0]  ( .D(\U4/Z_0 ), .CK(clock), .Q(\add_32/A[0] ), .QN(
        n549) );
  DFF_X1 \count_reg[1]  ( .D(\U4/Z_1 ), .CK(clock), .Q(\add_32/A[1] ), .QN(
        n548) );
  DFF_X1 \count_reg[2]  ( .D(\U4/Z_2 ), .CK(clock), .Q(\add_32/A[2] ) );
  DFF_X1 \count_reg[3]  ( .D(\U4/Z_3 ), .CK(clock), .Q(\add_32/A[3] ) );
  NOR2_X2 U99 ( .A1(\add_32/A[0] ), .A2(n29), .ZN(\U4/Z_0 ) );
  NOR2_X2 U101 ( .A1(set_bit), .A2(reset), .ZN(n32) );
  NAND4_X2 U102 ( .A1(n33), .A2(n34), .A3(n35), .A4(n36), .ZN(n31) );
  NOR3_X2 U103 ( .A1(element[18]), .A2(element[1]), .A3(element[19]), .ZN(n36)
         );
  NOR3_X2 U104 ( .A1(element[15]), .A2(element[17]), .A3(element[16]), .ZN(n35) );
  NOR3_X2 U105 ( .A1(element[12]), .A2(element[14]), .A3(element[13]), .ZN(n34) );
  NOR3_X2 U106 ( .A1(element[0]), .A2(element[11]), .A3(element[10]), .ZN(n33)
         );
  NAND4_X2 U107 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(n30) );
  NOR4_X2 U108 ( .A1(element[9]), .A2(element[8]), .A3(element[7]), .A4(
        element[6]), .ZN(n40) );
  NOR3_X2 U109 ( .A1(element[3]), .A2(element[5]), .A3(element[4]), .ZN(n39)
         );
  NOR3_X2 U110 ( .A1(element[23]), .A2(element[2]), .A3(element[24]), .ZN(n38)
         );
  NOR3_X2 U111 ( .A1(element[20]), .A2(element[22]), .A3(element[21]), .ZN(n37) );
  NOR2_X2 U112 ( .A1(n41), .A2(n567), .ZN(\U10/Z_9 ) );
  NOR2_X2 U113 ( .A1(n41), .A2(n568), .ZN(\U10/Z_8 ) );
  NOR2_X2 U114 ( .A1(n41), .A2(n569), .ZN(\U10/Z_7 ) );
  NOR2_X2 U115 ( .A1(n41), .A2(n570), .ZN(\U10/Z_6 ) );
  NOR2_X2 U116 ( .A1(n41), .A2(n571), .ZN(\U10/Z_5 ) );
  NOR2_X2 U117 ( .A1(n41), .A2(n572), .ZN(\U10/Z_4 ) );
  NOR2_X2 U118 ( .A1(n41), .A2(n573), .ZN(\U10/Z_3 ) );
  NOR2_X2 U119 ( .A1(n41), .A2(n553), .ZN(\U10/Z_23 ) );
  NOR2_X2 U120 ( .A1(n41), .A2(n554), .ZN(\U10/Z_22 ) );
  NOR2_X2 U121 ( .A1(n41), .A2(n555), .ZN(\U10/Z_21 ) );
  NOR2_X2 U122 ( .A1(n41), .A2(n556), .ZN(\U10/Z_20 ) );
  NOR2_X2 U123 ( .A1(n41), .A2(n574), .ZN(\U10/Z_2 ) );
  NOR2_X2 U124 ( .A1(n41), .A2(n557), .ZN(\U10/Z_19 ) );
  NOR2_X2 U125 ( .A1(n41), .A2(n558), .ZN(\U10/Z_18 ) );
  NOR2_X2 U126 ( .A1(n41), .A2(n559), .ZN(\U10/Z_17 ) );
  NOR2_X2 U127 ( .A1(n41), .A2(n560), .ZN(\U10/Z_16 ) );
  NOR2_X2 U128 ( .A1(n41), .A2(n561), .ZN(\U10/Z_15 ) );
  NOR2_X2 U129 ( .A1(n41), .A2(n562), .ZN(\U10/Z_14 ) );
  NOR2_X2 U130 ( .A1(n41), .A2(n563), .ZN(\U10/Z_13 ) );
  NOR2_X2 U131 ( .A1(n41), .A2(n564), .ZN(\U10/Z_12 ) );
  NOR2_X2 U132 ( .A1(n41), .A2(n565), .ZN(\U10/Z_11 ) );
  NOR2_X2 U133 ( .A1(n41), .A2(n566), .ZN(\U10/Z_10 ) );
  NOR2_X2 U134 ( .A1(n41), .A2(n575), .ZN(\U10/Z_1 ) );
  NOR2_X2 U135 ( .A1(n41), .A2(n576), .ZN(\U10/Z_0 ) );
  NAND2_X2 U136 ( .A1(n42), .A2(n552), .ZN(n41) );
  OAI33_X1 U164 ( .A1(n1), .A2(\add_32/carry[4] ), .A3(n29), .B1(n550), .B2(
        \add_32/A[4] ), .B3(n29), .ZN(n44) );
  AND2_X1 U165 ( .A1(\U4/DATA2_3 ), .A2(n551), .ZN(\U4/Z_3 ) );
  AND2_X1 U166 ( .A1(\U4/DATA2_2 ), .A2(n551), .ZN(\U4/Z_2 ) );
  AND2_X1 U167 ( .A1(\U4/DATA2_1 ), .A2(n551), .ZN(\U4/Z_1 ) );
  OR4_X1 U168 ( .A1(\add_32/A[2] ), .A2(n43), .A3(\add_32/A[4] ), .A4(
        \add_32/A[3] ), .ZN(n42) );
  DFF_X2 \count_reg[4]  ( .D(n44), .CK(clock), .Q(\add_32/A[4] ), .QN(n1) );
  INV_X4 U100 ( .A(1'b1), .ZN(adder_out4[0]) );
  INV_X4 U138 ( .A(1'b1), .ZN(adder_out4[1]) );
  INV_X4 U140 ( .A(1'b1), .ZN(adder_out4[2]) );
  INV_X4 U142 ( .A(1'b1), .ZN(adder_out4[3]) );
  INV_X4 U144 ( .A(1'b1), .ZN(adder_out4[4]) );
  INV_X4 U146 ( .A(1'b1), .ZN(adder_out4[5]) );
  INV_X4 U148 ( .A(1'b1), .ZN(adder_out4[6]) );
  INV_X4 U150 ( .A(1'b1), .ZN(adder_out4[7]) );
  INV_X4 U152 ( .A(1'b1), .ZN(adder_out4[8]) );
  INV_X4 U154 ( .A(1'b1), .ZN(adder_out4[9]) );
  INV_X4 U156 ( .A(1'b1), .ZN(adder_out4[10]) );
  INV_X4 U158 ( .A(1'b1), .ZN(adder_out4[11]) );
  INV_X4 U160 ( .A(1'b1), .ZN(adder_out4[12]) );
  INV_X4 U162 ( .A(1'b1), .ZN(adder_out4[13]) );
  INV_X4 U169 ( .A(1'b1), .ZN(adder_out4[14]) );
  INV_X4 U171 ( .A(1'b1), .ZN(adder_out4[15]) );
  INV_X4 U173 ( .A(1'b1), .ZN(adder_out4[16]) );
  INV_X4 U175 ( .A(1'b1), .ZN(adder_out4[17]) );
  INV_X4 U177 ( .A(1'b1), .ZN(adder_out4[18]) );
  INV_X4 U179 ( .A(1'b1), .ZN(adder_out4[19]) );
  INV_X4 U181 ( .A(1'b1), .ZN(adder_out4[20]) );
  INV_X4 U183 ( .A(1'b1), .ZN(adder_out4[21]) );
  INV_X4 U185 ( .A(1'b1), .ZN(adder_out4[22]) );
  INV_X4 U187 ( .A(1'b1), .ZN(adder_out4[23]) );
  INV_X4 U189 ( .A(1'b1), .ZN(adder_out3[0]) );
  INV_X4 U191 ( .A(1'b1), .ZN(adder_out3[1]) );
  INV_X4 U193 ( .A(1'b1), .ZN(adder_out3[2]) );
  INV_X4 U195 ( .A(1'b1), .ZN(adder_out3[3]) );
  INV_X4 U197 ( .A(1'b1), .ZN(adder_out3[4]) );
  INV_X4 U199 ( .A(1'b1), .ZN(adder_out3[5]) );
  INV_X4 U201 ( .A(1'b1), .ZN(adder_out3[6]) );
  INV_X4 U203 ( .A(1'b1), .ZN(adder_out3[7]) );
  INV_X4 U205 ( .A(1'b1), .ZN(adder_out3[8]) );
  INV_X4 U207 ( .A(1'b1), .ZN(adder_out3[9]) );
  INV_X4 U209 ( .A(1'b1), .ZN(adder_out3[10]) );
  INV_X4 U211 ( .A(1'b1), .ZN(adder_out3[11]) );
  INV_X4 U213 ( .A(1'b1), .ZN(adder_out3[12]) );
  INV_X4 U215 ( .A(1'b1), .ZN(adder_out3[13]) );
  INV_X4 U217 ( .A(1'b1), .ZN(adder_out3[14]) );
  INV_X4 U219 ( .A(1'b1), .ZN(adder_out3[15]) );
  INV_X4 U221 ( .A(1'b1), .ZN(adder_out3[16]) );
  INV_X4 U223 ( .A(1'b1), .ZN(adder_out3[17]) );
  INV_X4 U225 ( .A(1'b1), .ZN(adder_out3[18]) );
  INV_X4 U227 ( .A(1'b1), .ZN(adder_out3[19]) );
  INV_X4 U229 ( .A(1'b1), .ZN(adder_out3[20]) );
  INV_X4 U231 ( .A(1'b1), .ZN(adder_out3[21]) );
  INV_X4 U233 ( .A(1'b1), .ZN(adder_out3[22]) );
  INV_X4 U235 ( .A(1'b1), .ZN(adder_out3[23]) );
  INV_X4 U237 ( .A(1'b1), .ZN(adder_out2[0]) );
  INV_X4 U239 ( .A(1'b1), .ZN(adder_out2[1]) );
  INV_X4 U241 ( .A(1'b1), .ZN(adder_out2[2]) );
  INV_X4 U243 ( .A(1'b1), .ZN(adder_out2[3]) );
  INV_X4 U245 ( .A(1'b1), .ZN(adder_out2[4]) );
  INV_X4 U247 ( .A(1'b1), .ZN(adder_out2[5]) );
  INV_X4 U249 ( .A(1'b1), .ZN(adder_out2[6]) );
  INV_X4 U251 ( .A(1'b1), .ZN(adder_out2[7]) );
  INV_X4 U253 ( .A(1'b1), .ZN(adder_out2[8]) );
  INV_X4 U255 ( .A(1'b1), .ZN(adder_out2[9]) );
  INV_X4 U257 ( .A(1'b1), .ZN(adder_out2[10]) );
  INV_X4 U259 ( .A(1'b1), .ZN(adder_out2[11]) );
  INV_X4 U261 ( .A(1'b1), .ZN(adder_out2[12]) );
  INV_X4 U263 ( .A(1'b1), .ZN(adder_out2[13]) );
  INV_X4 U265 ( .A(1'b1), .ZN(adder_out2[14]) );
  INV_X4 U267 ( .A(1'b1), .ZN(adder_out2[15]) );
  INV_X4 U269 ( .A(1'b1), .ZN(adder_out2[16]) );
  INV_X4 U271 ( .A(1'b1), .ZN(adder_out2[17]) );
  INV_X4 U273 ( .A(1'b1), .ZN(adder_out2[18]) );
  INV_X4 U275 ( .A(1'b1), .ZN(adder_out2[19]) );
  INV_X4 U277 ( .A(1'b1), .ZN(adder_out2[20]) );
  INV_X4 U279 ( .A(1'b1), .ZN(adder_out2[21]) );
  INV_X4 U281 ( .A(1'b1), .ZN(adder_out2[22]) );
  INV_X4 U283 ( .A(1'b1), .ZN(adder_out2[23]) );
  INV_X4 U285 ( .A(1'b1), .ZN(adder_out1[0]) );
  INV_X4 U287 ( .A(1'b1), .ZN(adder_out1[1]) );
  INV_X4 U289 ( .A(1'b1), .ZN(adder_out1[2]) );
  INV_X4 U291 ( .A(1'b1), .ZN(adder_out1[3]) );
  INV_X4 U293 ( .A(1'b1), .ZN(adder_out1[4]) );
  INV_X4 U295 ( .A(1'b1), .ZN(adder_out1[5]) );
  INV_X4 U297 ( .A(1'b1), .ZN(adder_out1[6]) );
  INV_X4 U299 ( .A(1'b1), .ZN(adder_out1[7]) );
  INV_X4 U301 ( .A(1'b1), .ZN(adder_out1[8]) );
  INV_X4 U303 ( .A(1'b1), .ZN(adder_out1[9]) );
  INV_X4 U305 ( .A(1'b1), .ZN(adder_out1[10]) );
  INV_X4 U307 ( .A(1'b1), .ZN(adder_out1[11]) );
  INV_X4 U309 ( .A(1'b1), .ZN(adder_out1[12]) );
  INV_X4 U311 ( .A(1'b1), .ZN(adder_out1[13]) );
  INV_X4 U313 ( .A(1'b1), .ZN(adder_out1[14]) );
  INV_X4 U315 ( .A(1'b1), .ZN(adder_out1[15]) );
  INV_X4 U317 ( .A(1'b1), .ZN(adder_out1[16]) );
  INV_X4 U319 ( .A(1'b1), .ZN(adder_out1[17]) );
  INV_X4 U321 ( .A(1'b1), .ZN(adder_out1[18]) );
  INV_X4 U323 ( .A(1'b1), .ZN(adder_out1[19]) );
  INV_X4 U325 ( .A(1'b1), .ZN(adder_out1[20]) );
  INV_X4 U327 ( .A(1'b1), .ZN(adder_out1[21]) );
  INV_X4 U329 ( .A(1'b1), .ZN(adder_out1[22]) );
  INV_X4 U331 ( .A(1'b1), .ZN(adder_out1[23]) );
  NOR2_X2 U333 ( .A1(n548), .A2(n549), .ZN(n43) );
  OAI21_X2 U334 ( .B1(n30), .B2(n31), .A(n32), .ZN(n29) );
  INV_X4 U335 ( .A(\add_32/carry[4] ), .ZN(n550) );
  INV_X4 U336 ( .A(n29), .ZN(n551) );
  INV_X4 U337 ( .A(set_bit), .ZN(n552) );
  INV_X4 U338 ( .A(\U10/DATA2_23 ), .ZN(n553) );
  INV_X4 U339 ( .A(\U10/DATA2_22 ), .ZN(n554) );
  INV_X4 U340 ( .A(\U10/DATA2_21 ), .ZN(n555) );
  INV_X4 U341 ( .A(\U10/DATA2_20 ), .ZN(n556) );
  INV_X4 U342 ( .A(\U10/DATA2_19 ), .ZN(n557) );
  INV_X4 U343 ( .A(\U10/DATA2_18 ), .ZN(n558) );
  INV_X4 U344 ( .A(\U10/DATA2_17 ), .ZN(n559) );
  INV_X4 U345 ( .A(\U10/DATA2_16 ), .ZN(n560) );
  INV_X4 U346 ( .A(\U10/DATA2_15 ), .ZN(n561) );
  INV_X4 U347 ( .A(\U10/DATA2_14 ), .ZN(n562) );
  INV_X4 U348 ( .A(\U10/DATA2_13 ), .ZN(n563) );
  INV_X4 U349 ( .A(\U10/DATA2_12 ), .ZN(n564) );
  INV_X4 U350 ( .A(\U10/DATA2_11 ), .ZN(n565) );
  INV_X4 U351 ( .A(\U10/DATA2_10 ), .ZN(n566) );
  INV_X4 U352 ( .A(\U10/DATA2_9 ), .ZN(n567) );
  INV_X4 U353 ( .A(\U10/DATA2_8 ), .ZN(n568) );
  INV_X4 U354 ( .A(\U10/DATA2_7 ), .ZN(n569) );
  INV_X4 U355 ( .A(\U10/DATA2_6 ), .ZN(n570) );
  INV_X4 U356 ( .A(\U10/DATA2_5 ), .ZN(n571) );
  INV_X4 U357 ( .A(\U10/DATA2_4 ), .ZN(n572) );
  INV_X4 U358 ( .A(\U10/DATA2_3 ), .ZN(n573) );
  INV_X4 U359 ( .A(\U10/DATA2_2 ), .ZN(n574) );
  INV_X4 U360 ( .A(\U10/DATA2_1 ), .ZN(n575) );
  INV_X4 U361 ( .A(\U10/DATA2_0 ), .ZN(n576) );
endmodule


module syncAccum_1 ( clock, mult_output, accum_input, accum_output, 
        accum_output25 );
  input [24:0] mult_output;
  output [23:0] accum_input;
  input [23:0] accum_output;
  output [24:0] accum_output25;
  input clock;
  wire   dirtybuff1, dirtybuff2, dirtybuff3;

  DFF_X1 dirtybuff1_reg ( .D(mult_output[24]), .CK(clock), .Q(dirtybuff1) );
  DFF_X1 dirtybuff2_reg ( .D(dirtybuff1), .CK(clock), .Q(dirtybuff2) );
  DFF_X1 dirtybuff3_reg ( .D(dirtybuff2), .CK(clock), .Q(dirtybuff3) );
  DFF_X1 dirtybuff4_reg ( .D(dirtybuff3), .CK(clock), .Q(accum_output25[24])
         );
  BUF_X4 U3 ( .A(mult_output[0]), .Z(accum_input[0]) );
  BUF_X4 U4 ( .A(mult_output[1]), .Z(accum_input[1]) );
  BUF_X4 U5 ( .A(mult_output[2]), .Z(accum_input[2]) );
  BUF_X4 U6 ( .A(mult_output[3]), .Z(accum_input[3]) );
  BUF_X4 U7 ( .A(mult_output[4]), .Z(accum_input[4]) );
  BUF_X4 U8 ( .A(mult_output[5]), .Z(accum_input[5]) );
  BUF_X4 U9 ( .A(mult_output[6]), .Z(accum_input[6]) );
  BUF_X4 U10 ( .A(mult_output[7]), .Z(accum_input[7]) );
  BUF_X4 U11 ( .A(mult_output[8]), .Z(accum_input[8]) );
  BUF_X4 U12 ( .A(mult_output[9]), .Z(accum_input[9]) );
  BUF_X4 U13 ( .A(mult_output[10]), .Z(accum_input[10]) );
  BUF_X4 U14 ( .A(mult_output[11]), .Z(accum_input[11]) );
  BUF_X4 U15 ( .A(mult_output[12]), .Z(accum_input[12]) );
  BUF_X4 U16 ( .A(mult_output[13]), .Z(accum_input[13]) );
  BUF_X4 U17 ( .A(mult_output[14]), .Z(accum_input[14]) );
  BUF_X4 U18 ( .A(mult_output[15]), .Z(accum_input[15]) );
  BUF_X4 U19 ( .A(mult_output[16]), .Z(accum_input[16]) );
  BUF_X4 U20 ( .A(mult_output[17]), .Z(accum_input[17]) );
  BUF_X4 U21 ( .A(mult_output[18]), .Z(accum_input[18]) );
  BUF_X4 U22 ( .A(mult_output[19]), .Z(accum_input[19]) );
  BUF_X4 U23 ( .A(mult_output[20]), .Z(accum_input[20]) );
  BUF_X4 U24 ( .A(mult_output[21]), .Z(accum_input[21]) );
  BUF_X4 U25 ( .A(mult_output[22]), .Z(accum_input[22]) );
  BUF_X4 U26 ( .A(mult_output[23]), .Z(accum_input[23]) );
  BUF_X4 U27 ( .A(accum_output[0]), .Z(accum_output25[0]) );
  BUF_X4 U28 ( .A(accum_output[1]), .Z(accum_output25[1]) );
  BUF_X4 U29 ( .A(accum_output[2]), .Z(accum_output25[2]) );
  BUF_X4 U30 ( .A(accum_output[3]), .Z(accum_output25[3]) );
  BUF_X4 U31 ( .A(accum_output[4]), .Z(accum_output25[4]) );
  BUF_X4 U32 ( .A(accum_output[5]), .Z(accum_output25[5]) );
  BUF_X4 U33 ( .A(accum_output[6]), .Z(accum_output25[6]) );
  BUF_X4 U34 ( .A(accum_output[7]), .Z(accum_output25[7]) );
  BUF_X4 U35 ( .A(accum_output[8]), .Z(accum_output25[8]) );
  BUF_X4 U36 ( .A(accum_output[9]), .Z(accum_output25[9]) );
  BUF_X4 U37 ( .A(accum_output[10]), .Z(accum_output25[10]) );
  BUF_X4 U38 ( .A(accum_output[11]), .Z(accum_output25[11]) );
  BUF_X4 U39 ( .A(accum_output[12]), .Z(accum_output25[12]) );
  BUF_X4 U40 ( .A(accum_output[13]), .Z(accum_output25[13]) );
  BUF_X4 U41 ( .A(accum_output[14]), .Z(accum_output25[14]) );
  BUF_X4 U42 ( .A(accum_output[15]), .Z(accum_output25[15]) );
  BUF_X4 U43 ( .A(accum_output[16]), .Z(accum_output25[16]) );
  BUF_X4 U44 ( .A(accum_output[17]), .Z(accum_output25[17]) );
  BUF_X4 U45 ( .A(accum_output[18]), .Z(accum_output25[18]) );
  BUF_X4 U46 ( .A(accum_output[19]), .Z(accum_output25[19]) );
  BUF_X4 U47 ( .A(accum_output[20]), .Z(accum_output25[20]) );
  BUF_X4 U48 ( .A(accum_output[21]), .Z(accum_output25[21]) );
  BUF_X4 U49 ( .A(accum_output[22]), .Z(accum_output25[22]) );
  BUF_X4 U50 ( .A(accum_output[23]), .Z(accum_output25[23]) );
endmodule


module isched ( clock, reset, addressI, data, dataI, FinalOutput, sig );
  output [7:0] addressI;
  input [191:0] data;
  output [47:0] dataI;
  input [23:0] FinalOutput;
  input clock, reset, sig;
  wire   n96, \U13/DATA2_0 , \U7/Z_0 , \U7/Z_1 , \U7/Z_2 , \U7/Z_3 , \U7/Z_4 ,
         \U7/Z_5 , \U7/Z_6 , \U7/Z_7 , \U7/Z_8 , \U7/Z_9 , \U7/Z_10 ,
         \U7/Z_11 , \U7/Z_12 , \U7/Z_13 , \U7/Z_14 , \U7/Z_15 , \U7/Z_16 ,
         \U7/Z_17 , \U7/Z_18 , \U7/Z_19 , \U7/Z_20 , \U7/Z_21 , \U7/Z_22 ,
         \U7/Z_23 , \U7/Z_24 , \U7/Z_25 , \U7/Z_26 , \U7/Z_27 , \U7/Z_28 ,
         \U7/Z_29 , \U7/Z_30 , \U7/Z_31 , \U7/Z_32 , \U7/Z_33 , \U7/Z_34 ,
         \U7/Z_35 , \U7/Z_36 , \U7/Z_37 , \U7/Z_38 , \U7/Z_39 , \U7/Z_40 ,
         \U7/Z_41 , \U7/Z_42 , \U7/Z_43 , \U7/Z_44 , \U7/Z_45 , \U7/Z_46 ,
         \U7/Z_47 , \U7/DATA5_0 , \U7/DATA5_1 , \U7/DATA5_2 , \U7/DATA5_3 ,
         \U7/DATA5_4 , \U7/DATA5_5 , \U7/DATA5_6 , \U7/DATA5_7 , \U7/DATA5_8 ,
         \U7/DATA5_9 , \U7/DATA5_10 , \U7/DATA5_11 , \U7/DATA5_12 ,
         \U7/DATA5_13 , \U7/DATA5_14 , \U7/DATA5_15 , \U7/DATA5_16 ,
         \U7/DATA5_17 , \U7/DATA5_18 , \U7/DATA5_19 , \U7/DATA5_20 ,
         \U7/DATA5_21 , \U7/DATA5_22 , \U7/DATA5_23 , \U7/DATA5_24 ,
         \U7/DATA5_25 , \U7/DATA5_26 , \U7/DATA5_27 , \U7/DATA5_28 ,
         \U7/DATA5_29 , \U7/DATA5_30 , \U7/DATA5_31 , \U7/DATA5_32 ,
         \U7/DATA5_33 , \U7/DATA5_34 , \U7/DATA5_35 , \U7/DATA5_36 ,
         \U7/DATA5_37 , \U7/DATA5_38 , \U7/DATA5_39 , \U7/DATA5_40 ,
         \U7/DATA5_41 , \U7/DATA5_42 , \U7/DATA5_43 , \U7/DATA5_44 ,
         \U7/DATA5_45 , \U7/DATA5_46 , \U7/DATA5_47 , \U7/DATA4_0 ,
         \U7/DATA4_1 , \U7/DATA4_2 , \U7/DATA4_3 , \U7/DATA4_4 , \U7/DATA4_5 ,
         \U7/DATA4_6 , \U7/DATA4_7 , \U7/DATA4_8 , \U7/DATA4_9 , \U7/DATA4_10 ,
         \U7/DATA4_11 , \U7/DATA4_12 , \U7/DATA4_13 , \U7/DATA4_14 ,
         \U7/DATA4_15 , \U7/DATA4_16 , \U7/DATA4_17 , \U7/DATA4_18 ,
         \U7/DATA4_19 , \U7/DATA4_20 , \U7/DATA4_21 , \U7/DATA4_22 ,
         \U7/DATA4_23 , \U7/DATA4_24 , \U7/DATA4_25 , \U7/DATA4_26 ,
         \U7/DATA4_27 , \U7/DATA4_28 , \U7/DATA4_29 , \U7/DATA4_30 ,
         \U7/DATA4_31 , \U7/DATA4_32 , \U7/DATA4_33 , \U7/DATA4_34 ,
         \U7/DATA4_35 , \U7/DATA4_36 , \U7/DATA4_37 , \U7/DATA4_38 ,
         \U7/DATA4_39 , \U7/DATA4_40 , \U7/DATA4_41 , \U7/DATA4_42 ,
         \U7/DATA4_43 , \U7/DATA4_44 , \U7/DATA4_45 , \U7/DATA4_46 ,
         \U7/DATA4_47 , \U7/DATA3_0 , \U7/DATA3_1 , \U7/DATA3_2 , \U7/DATA3_3 ,
         \U7/DATA3_4 , \U7/DATA3_5 , \U7/DATA3_6 , \U7/DATA3_7 , \U7/DATA3_8 ,
         \U7/DATA3_9 , \U7/DATA3_10 , \U7/DATA3_11 , \U7/DATA3_12 ,
         \U7/DATA3_13 , \U7/DATA3_14 , \U7/DATA3_15 , \U7/DATA3_16 ,
         \U7/DATA3_17 , \U7/DATA3_18 , \U7/DATA3_19 , \U7/DATA3_20 ,
         \U7/DATA3_21 , \U7/DATA3_22 , \U7/DATA3_23 , \U7/DATA3_24 ,
         \U7/DATA3_25 , \U7/DATA3_26 , \U7/DATA3_27 , \U7/DATA3_28 ,
         \U7/DATA3_29 , \U7/DATA3_30 , \U7/DATA3_31 , \U7/DATA3_32 ,
         \U7/DATA3_33 , \U7/DATA3_34 , \U7/DATA3_35 , \U7/DATA3_36 ,
         \U7/DATA3_37 , \U7/DATA3_38 , \U7/DATA3_39 , \U7/DATA3_40 ,
         \U7/DATA3_41 , \U7/DATA3_42 , \U7/DATA3_43 , \U7/DATA3_44 ,
         \U7/DATA3_45 , \U7/DATA3_46 , \U7/DATA3_47 , \U7/DATA2_0 ,
         \U7/DATA2_1 , \U7/DATA2_2 , \U7/DATA2_3 , \U7/DATA2_4 , \U7/DATA2_5 ,
         \U7/DATA2_6 , \U7/DATA2_7 , \U7/DATA2_8 , \U7/DATA2_9 , \U7/DATA2_10 ,
         \U7/DATA2_11 , \U7/DATA2_12 , \U7/DATA2_13 , \U7/DATA2_14 ,
         \U7/DATA2_15 , \U7/DATA2_16 , \U7/DATA2_17 , \U7/DATA2_18 ,
         \U7/DATA2_19 , \U7/DATA2_20 , \U7/DATA2_21 , \U7/DATA2_22 ,
         \U7/DATA2_23 , \U7/DATA2_24 , \U7/DATA2_25 , \U7/DATA2_26 ,
         \U7/DATA2_27 , \U7/DATA2_28 , \U7/DATA2_29 , \U7/DATA2_30 ,
         \U7/DATA2_31 , \U7/DATA2_32 , \U7/DATA2_33 , \U7/DATA2_34 ,
         \U7/DATA2_35 , \U7/DATA2_36 , \U7/DATA2_37 , \U7/DATA2_38 ,
         \U7/DATA2_39 , \U7/DATA2_40 , \U7/DATA2_41 , \U7/DATA2_42 ,
         \U7/DATA2_43 , \U7/DATA2_44 , \U7/DATA2_45 , \U7/DATA2_46 ,
         \U7/DATA2_47 , \U4/DATA1_1 , \U4/DATA1_2 , \U4/DATA1_3 , \U4/DATA1_4 ,
         \U4/DATA1_5 , \U4/DATA1_6 , \add_54/carry[7] , \add_54/carry[6] ,
         \add_54/carry[5] , \add_54/carry[4] , \add_54/carry[3] ,
         \add_54/carry[2] , \add_54/A[0] , \add_54/A[1] , \add_54/A[2] ,
         \add_54/A[3] , \add_54/A[4] , \add_54/A[5] , \add_54/A[6] ,
         \add_54/A[7] , \add_46/A[0] , \add_46/A[1] , \add_46/A[2] , n12, n13,
         n15, n16, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n55, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402;
  assign \U13/DATA2_0  = reset;
  assign dataI[0] = \U7/Z_0 ;
  assign dataI[1] = \U7/Z_1 ;
  assign dataI[2] = \U7/Z_2 ;
  assign dataI[3] = \U7/Z_3 ;
  assign dataI[4] = \U7/Z_4 ;
  assign dataI[5] = \U7/Z_5 ;
  assign dataI[6] = \U7/Z_6 ;
  assign dataI[7] = \U7/Z_7 ;
  assign dataI[8] = \U7/Z_8 ;
  assign dataI[9] = \U7/Z_9 ;
  assign dataI[10] = \U7/Z_10 ;
  assign dataI[11] = \U7/Z_11 ;
  assign dataI[12] = \U7/Z_12 ;
  assign dataI[13] = \U7/Z_13 ;
  assign dataI[14] = \U7/Z_14 ;
  assign dataI[15] = \U7/Z_15 ;
  assign dataI[16] = \U7/Z_16 ;
  assign dataI[17] = \U7/Z_17 ;
  assign dataI[18] = \U7/Z_18 ;
  assign dataI[19] = \U7/Z_19 ;
  assign dataI[20] = \U7/Z_20 ;
  assign dataI[21] = \U7/Z_21 ;
  assign dataI[22] = \U7/Z_22 ;
  assign dataI[23] = \U7/Z_23 ;
  assign dataI[24] = \U7/Z_24 ;
  assign dataI[25] = \U7/Z_25 ;
  assign dataI[26] = \U7/Z_26 ;
  assign dataI[27] = \U7/Z_27 ;
  assign dataI[28] = \U7/Z_28 ;
  assign dataI[29] = \U7/Z_29 ;
  assign dataI[30] = \U7/Z_30 ;
  assign dataI[31] = \U7/Z_31 ;
  assign dataI[32] = \U7/Z_32 ;
  assign dataI[33] = \U7/Z_33 ;
  assign dataI[34] = \U7/Z_34 ;
  assign dataI[35] = \U7/Z_35 ;
  assign dataI[36] = \U7/Z_36 ;
  assign dataI[37] = \U7/Z_37 ;
  assign dataI[38] = \U7/Z_38 ;
  assign dataI[39] = \U7/Z_39 ;
  assign dataI[40] = \U7/Z_40 ;
  assign dataI[41] = \U7/Z_41 ;
  assign dataI[42] = \U7/Z_42 ;
  assign dataI[43] = \U7/Z_43 ;
  assign dataI[44] = \U7/Z_44 ;
  assign dataI[45] = \U7/Z_45 ;
  assign dataI[46] = \U7/Z_46 ;
  assign dataI[47] = \U7/Z_47 ;
  assign \U7/DATA5_0  = data[0];
  assign \U7/DATA5_1  = data[1];
  assign \U7/DATA5_2  = data[2];
  assign \U7/DATA5_3  = data[3];
  assign \U7/DATA5_4  = data[4];
  assign \U7/DATA5_5  = data[5];
  assign \U7/DATA5_6  = data[6];
  assign \U7/DATA5_7  = data[7];
  assign \U7/DATA5_8  = data[8];
  assign \U7/DATA5_9  = data[9];
  assign \U7/DATA5_10  = data[10];
  assign \U7/DATA5_11  = data[11];
  assign \U7/DATA5_12  = data[12];
  assign \U7/DATA5_13  = data[13];
  assign \U7/DATA5_14  = data[14];
  assign \U7/DATA5_15  = data[15];
  assign \U7/DATA5_16  = data[16];
  assign \U7/DATA5_17  = data[17];
  assign \U7/DATA5_18  = data[18];
  assign \U7/DATA5_19  = data[19];
  assign \U7/DATA5_20  = data[20];
  assign \U7/DATA5_21  = data[21];
  assign \U7/DATA5_22  = data[22];
  assign \U7/DATA5_23  = data[23];
  assign \U7/DATA5_24  = data[24];
  assign \U7/DATA5_25  = data[25];
  assign \U7/DATA5_26  = data[26];
  assign \U7/DATA5_27  = data[27];
  assign \U7/DATA5_28  = data[28];
  assign \U7/DATA5_29  = data[29];
  assign \U7/DATA5_30  = data[30];
  assign \U7/DATA5_31  = data[31];
  assign \U7/DATA5_32  = data[32];
  assign \U7/DATA5_33  = data[33];
  assign \U7/DATA5_34  = data[34];
  assign \U7/DATA5_35  = data[35];
  assign \U7/DATA5_36  = data[36];
  assign \U7/DATA5_37  = data[37];
  assign \U7/DATA5_38  = data[38];
  assign \U7/DATA5_39  = data[39];
  assign \U7/DATA5_40  = data[40];
  assign \U7/DATA5_41  = data[41];
  assign \U7/DATA5_42  = data[42];
  assign \U7/DATA5_43  = data[43];
  assign \U7/DATA5_44  = data[44];
  assign \U7/DATA5_45  = data[45];
  assign \U7/DATA5_46  = data[46];
  assign \U7/DATA5_47  = data[47];
  assign \U7/DATA4_0  = data[48];
  assign \U7/DATA4_1  = data[49];
  assign \U7/DATA4_2  = data[50];
  assign \U7/DATA4_3  = data[51];
  assign \U7/DATA4_4  = data[52];
  assign \U7/DATA4_5  = data[53];
  assign \U7/DATA4_6  = data[54];
  assign \U7/DATA4_7  = data[55];
  assign \U7/DATA4_8  = data[56];
  assign \U7/DATA4_9  = data[57];
  assign \U7/DATA4_10  = data[58];
  assign \U7/DATA4_11  = data[59];
  assign \U7/DATA4_12  = data[60];
  assign \U7/DATA4_13  = data[61];
  assign \U7/DATA4_14  = data[62];
  assign \U7/DATA4_15  = data[63];
  assign \U7/DATA4_16  = data[64];
  assign \U7/DATA4_17  = data[65];
  assign \U7/DATA4_18  = data[66];
  assign \U7/DATA4_19  = data[67];
  assign \U7/DATA4_20  = data[68];
  assign \U7/DATA4_21  = data[69];
  assign \U7/DATA4_22  = data[70];
  assign \U7/DATA4_23  = data[71];
  assign \U7/DATA4_24  = data[72];
  assign \U7/DATA4_25  = data[73];
  assign \U7/DATA4_26  = data[74];
  assign \U7/DATA4_27  = data[75];
  assign \U7/DATA4_28  = data[76];
  assign \U7/DATA4_29  = data[77];
  assign \U7/DATA4_30  = data[78];
  assign \U7/DATA4_31  = data[79];
  assign \U7/DATA4_32  = data[80];
  assign \U7/DATA4_33  = data[81];
  assign \U7/DATA4_34  = data[82];
  assign \U7/DATA4_35  = data[83];
  assign \U7/DATA4_36  = data[84];
  assign \U7/DATA4_37  = data[85];
  assign \U7/DATA4_38  = data[86];
  assign \U7/DATA4_39  = data[87];
  assign \U7/DATA4_40  = data[88];
  assign \U7/DATA4_41  = data[89];
  assign \U7/DATA4_42  = data[90];
  assign \U7/DATA4_43  = data[91];
  assign \U7/DATA4_44  = data[92];
  assign \U7/DATA4_45  = data[93];
  assign \U7/DATA4_46  = data[94];
  assign \U7/DATA4_47  = data[95];
  assign \U7/DATA3_0  = data[96];
  assign \U7/DATA3_1  = data[97];
  assign \U7/DATA3_2  = data[98];
  assign \U7/DATA3_3  = data[99];
  assign \U7/DATA3_4  = data[100];
  assign \U7/DATA3_5  = data[101];
  assign \U7/DATA3_6  = data[102];
  assign \U7/DATA3_7  = data[103];
  assign \U7/DATA3_8  = data[104];
  assign \U7/DATA3_9  = data[105];
  assign \U7/DATA3_10  = data[106];
  assign \U7/DATA3_11  = data[107];
  assign \U7/DATA3_12  = data[108];
  assign \U7/DATA3_13  = data[109];
  assign \U7/DATA3_14  = data[110];
  assign \U7/DATA3_15  = data[111];
  assign \U7/DATA3_16  = data[112];
  assign \U7/DATA3_17  = data[113];
  assign \U7/DATA3_18  = data[114];
  assign \U7/DATA3_19  = data[115];
  assign \U7/DATA3_20  = data[116];
  assign \U7/DATA3_21  = data[117];
  assign \U7/DATA3_22  = data[118];
  assign \U7/DATA3_23  = data[119];
  assign \U7/DATA3_24  = data[120];
  assign \U7/DATA3_25  = data[121];
  assign \U7/DATA3_26  = data[122];
  assign \U7/DATA3_27  = data[123];
  assign \U7/DATA3_28  = data[124];
  assign \U7/DATA3_29  = data[125];
  assign \U7/DATA3_30  = data[126];
  assign \U7/DATA3_31  = data[127];
  assign \U7/DATA3_32  = data[128];
  assign \U7/DATA3_33  = data[129];
  assign \U7/DATA3_34  = data[130];
  assign \U7/DATA3_35  = data[131];
  assign \U7/DATA3_36  = data[132];
  assign \U7/DATA3_37  = data[133];
  assign \U7/DATA3_38  = data[134];
  assign \U7/DATA3_39  = data[135];
  assign \U7/DATA3_40  = data[136];
  assign \U7/DATA3_41  = data[137];
  assign \U7/DATA3_42  = data[138];
  assign \U7/DATA3_43  = data[139];
  assign \U7/DATA3_44  = data[140];
  assign \U7/DATA3_45  = data[141];
  assign \U7/DATA3_46  = data[142];
  assign \U7/DATA3_47  = data[143];
  assign \U7/DATA2_0  = data[144];
  assign \U7/DATA2_1  = data[145];
  assign \U7/DATA2_2  = data[146];
  assign \U7/DATA2_3  = data[147];
  assign \U7/DATA2_4  = data[148];
  assign \U7/DATA2_5  = data[149];
  assign \U7/DATA2_6  = data[150];
  assign \U7/DATA2_7  = data[151];
  assign \U7/DATA2_8  = data[152];
  assign \U7/DATA2_9  = data[153];
  assign \U7/DATA2_10  = data[154];
  assign \U7/DATA2_11  = data[155];
  assign \U7/DATA2_12  = data[156];
  assign \U7/DATA2_13  = data[157];
  assign \U7/DATA2_14  = data[158];
  assign \U7/DATA2_15  = data[159];
  assign \U7/DATA2_16  = data[160];
  assign \U7/DATA2_17  = data[161];
  assign \U7/DATA2_18  = data[162];
  assign \U7/DATA2_19  = data[163];
  assign \U7/DATA2_20  = data[164];
  assign \U7/DATA2_21  = data[165];
  assign \U7/DATA2_22  = data[166];
  assign \U7/DATA2_23  = data[167];
  assign \U7/DATA2_24  = data[168];
  assign \U7/DATA2_25  = data[169];
  assign \U7/DATA2_26  = data[170];
  assign \U7/DATA2_27  = data[171];
  assign \U7/DATA2_28  = data[172];
  assign \U7/DATA2_29  = data[173];
  assign \U7/DATA2_30  = data[174];
  assign \U7/DATA2_31  = data[175];
  assign \U7/DATA2_32  = data[176];
  assign \U7/DATA2_33  = data[177];
  assign \U7/DATA2_34  = data[178];
  assign \U7/DATA2_35  = data[179];
  assign \U7/DATA2_36  = data[180];
  assign \U7/DATA2_37  = data[181];
  assign \U7/DATA2_38  = data[182];
  assign \U7/DATA2_39  = data[183];
  assign \U7/DATA2_40  = data[184];
  assign \U7/DATA2_41  = data[185];
  assign \U7/DATA2_42  = data[186];
  assign \U7/DATA2_43  = data[187];
  assign \U7/DATA2_44  = data[188];
  assign \U7/DATA2_45  = data[189];
  assign \U7/DATA2_46  = data[190];
  assign \U7/DATA2_47  = data[191];
  assign addressI[0] = \add_54/A[0] ;
  assign addressI[1] = \add_54/A[1] ;
  assign addressI[2] = \add_54/A[2] ;
  assign addressI[3] = \add_54/A[3] ;
  assign addressI[4] = \add_54/A[4] ;
  assign addressI[5] = \add_54/A[5] ;
  assign addressI[6] = \add_54/A[6] ;
  assign addressI[7] = \add_54/A[7] ;

  HA_X1 \add_54/U1_1_1  ( .A(\add_54/A[1] ), .B(\add_54/A[0] ), .CO(
        \add_54/carry[2] ), .S(\U4/DATA1_1 ) );
  HA_X1 \add_54/U1_1_2  ( .A(\add_54/A[2] ), .B(\add_54/carry[2] ), .CO(
        \add_54/carry[3] ), .S(\U4/DATA1_2 ) );
  HA_X1 \add_54/U1_1_3  ( .A(\add_54/A[3] ), .B(\add_54/carry[3] ), .CO(
        \add_54/carry[4] ), .S(\U4/DATA1_3 ) );
  HA_X1 \add_54/U1_1_4  ( .A(\add_54/A[4] ), .B(\add_54/carry[4] ), .CO(
        \add_54/carry[5] ), .S(\U4/DATA1_4 ) );
  HA_X1 \add_54/U1_1_5  ( .A(\add_54/A[5] ), .B(\add_54/carry[5] ), .CO(
        \add_54/carry[6] ), .S(\U4/DATA1_5 ) );
  HA_X1 \add_54/U1_1_6  ( .A(\add_54/A[6] ), .B(\add_54/carry[6] ), .CO(
        \add_54/carry[7] ), .S(\U4/DATA1_6 ) );
  DFF_X2 NewRowFlag_reg ( .D(n157), .CK(clock), .Q(n384), .QN(n16) );
  DFF_X1 FirstFlag_reg ( .D(n158), .CK(clock), .Q(n96), .QN(n18) );
  DFF_X1 \count_reg[2]  ( .D(n156), .CK(clock), .Q(\add_46/A[2] ), .QN(n12) );
  DFF_X1 \count_reg[0]  ( .D(n154), .CK(clock), .Q(\add_46/A[0] ), .QN(n15) );
  DFF_X1 \count_reg[1]  ( .D(n155), .CK(clock), .Q(\add_46/A[1] ), .QN(n13) );
  NAND3_X2 U4 ( .A1(n23), .A2(n19), .A3(\add_54/carry[7] ), .ZN(n22) );
  OAI22_X2 U12 ( .A1(n390), .A2(n20), .B1(\add_54/A[0] ), .B2(n401), .ZN(n153)
         );
  NOR2_X2 U13 ( .A1(n398), .A2(n23), .ZN(n26) );
  OAI22_X2 U14 ( .A1(n32), .A2(n15), .B1(n23), .B2(n399), .ZN(n154) );
  NAND3_X2 U17 ( .A1(\add_46/A[0] ), .A2(n13), .A3(n37), .ZN(n36) );
  OAI22_X2 U18 ( .A1(n39), .A2(n12), .B1(n400), .B2(n40), .ZN(n156) );
  NAND3_X2 U21 ( .A1(n401), .A2(n34), .A3(n41), .ZN(n32) );
  NOR3_X2 U22 ( .A1(n398), .A2(sig), .A3(\U13/DATA2_0 ), .ZN(n41) );
  NOR2_X2 U23 ( .A1(n34), .A2(n23), .ZN(n37) );
  NAND3_X2 U24 ( .A1(n157), .A2(n402), .A3(n96), .ZN(n34) );
  NAND2_X2 U25 ( .A1(n42), .A2(n35), .ZN(n158) );
  NAND3_X2 U26 ( .A1(n18), .A2(n402), .A3(n157), .ZN(n35) );
  NAND4_X2 U27 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(n157) );
  NOR4_X2 U28 ( .A1(n47), .A2(FinalOutput[4]), .A3(FinalOutput[6]), .A4(
        FinalOutput[5]), .ZN(n46) );
  NOR4_X2 U29 ( .A1(n48), .A2(FinalOutput[20]), .A3(FinalOutput[22]), .A4(
        FinalOutput[21]), .ZN(n45) );
  NOR4_X2 U30 ( .A1(n49), .A2(FinalOutput[15]), .A3(FinalOutput[17]), .A4(
        FinalOutput[16]), .ZN(n44) );
  NOR4_X2 U31 ( .A1(n50), .A2(FinalOutput[0]), .A3(FinalOutput[11]), .A4(
        FinalOutput[10]), .ZN(n43) );
  NAND2_X2 U32 ( .A1(n51), .A2(n52), .ZN(\U7/Z_9 ) );
  NAND2_X2 U35 ( .A1(n57), .A2(n58), .ZN(\U7/Z_8 ) );
  NAND2_X2 U38 ( .A1(n59), .A2(n60), .ZN(\U7/Z_7 ) );
  NAND2_X2 U41 ( .A1(n61), .A2(n62), .ZN(\U7/Z_6 ) );
  NAND2_X2 U44 ( .A1(n63), .A2(n64), .ZN(\U7/Z_5 ) );
  NAND2_X2 U47 ( .A1(n65), .A2(n66), .ZN(\U7/Z_47 ) );
  NAND2_X2 U50 ( .A1(n67), .A2(n68), .ZN(\U7/Z_46 ) );
  NAND2_X2 U53 ( .A1(n69), .A2(n70), .ZN(\U7/Z_45 ) );
  NAND2_X2 U56 ( .A1(n71), .A2(n72), .ZN(\U7/Z_44 ) );
  NAND2_X2 U59 ( .A1(n73), .A2(n74), .ZN(\U7/Z_43 ) );
  NAND2_X2 U62 ( .A1(n75), .A2(n76), .ZN(\U7/Z_42 ) );
  NAND2_X2 U65 ( .A1(n77), .A2(n78), .ZN(\U7/Z_41 ) );
  NAND2_X2 U68 ( .A1(n79), .A2(n80), .ZN(\U7/Z_40 ) );
  NAND2_X2 U71 ( .A1(n81), .A2(n82), .ZN(\U7/Z_4 ) );
  NAND2_X2 U74 ( .A1(n83), .A2(n84), .ZN(\U7/Z_39 ) );
  NAND2_X2 U77 ( .A1(n85), .A2(n86), .ZN(\U7/Z_38 ) );
  NAND2_X2 U80 ( .A1(n87), .A2(n88), .ZN(\U7/Z_37 ) );
  NAND2_X2 U83 ( .A1(n89), .A2(n90), .ZN(\U7/Z_36 ) );
  NAND2_X2 U86 ( .A1(n91), .A2(n92), .ZN(\U7/Z_35 ) );
  NAND2_X2 U89 ( .A1(n93), .A2(n94), .ZN(\U7/Z_34 ) );
  NAND2_X2 U92 ( .A1(n95), .A2(n97), .ZN(\U7/Z_33 ) );
  NAND2_X2 U95 ( .A1(n98), .A2(n99), .ZN(\U7/Z_32 ) );
  NAND2_X2 U98 ( .A1(n100), .A2(n101), .ZN(\U7/Z_31 ) );
  NAND2_X2 U101 ( .A1(n102), .A2(n103), .ZN(\U7/Z_30 ) );
  NAND2_X2 U104 ( .A1(n104), .A2(n105), .ZN(\U7/Z_3 ) );
  NAND2_X2 U107 ( .A1(n106), .A2(n107), .ZN(\U7/Z_29 ) );
  NAND2_X2 U110 ( .A1(n108), .A2(n109), .ZN(\U7/Z_28 ) );
  NAND2_X2 U113 ( .A1(n110), .A2(n111), .ZN(\U7/Z_27 ) );
  NAND2_X2 U116 ( .A1(n112), .A2(n113), .ZN(\U7/Z_26 ) );
  NAND2_X2 U119 ( .A1(n114), .A2(n115), .ZN(\U7/Z_25 ) );
  NAND2_X2 U122 ( .A1(n116), .A2(n117), .ZN(\U7/Z_24 ) );
  NAND2_X2 U125 ( .A1(n118), .A2(n119), .ZN(\U7/Z_23 ) );
  NAND2_X2 U128 ( .A1(n120), .A2(n121), .ZN(\U7/Z_22 ) );
  NAND2_X2 U131 ( .A1(n122), .A2(n123), .ZN(\U7/Z_21 ) );
  NAND2_X2 U134 ( .A1(n124), .A2(n125), .ZN(\U7/Z_20 ) );
  NAND2_X2 U137 ( .A1(n126), .A2(n127), .ZN(\U7/Z_2 ) );
  NAND2_X2 U140 ( .A1(n128), .A2(n129), .ZN(\U7/Z_19 ) );
  NAND2_X2 U143 ( .A1(n130), .A2(n131), .ZN(\U7/Z_18 ) );
  NAND2_X2 U146 ( .A1(n132), .A2(n133), .ZN(\U7/Z_17 ) );
  NAND2_X2 U149 ( .A1(n134), .A2(n135), .ZN(\U7/Z_16 ) );
  NAND2_X2 U152 ( .A1(n136), .A2(n137), .ZN(\U7/Z_15 ) );
  NAND2_X2 U155 ( .A1(n138), .A2(n139), .ZN(\U7/Z_14 ) );
  NAND2_X2 U158 ( .A1(n140), .A2(n141), .ZN(\U7/Z_13 ) );
  NAND2_X2 U161 ( .A1(n142), .A2(n143), .ZN(\U7/Z_12 ) );
  NAND2_X2 U164 ( .A1(n144), .A2(n145), .ZN(\U7/Z_11 ) );
  NAND2_X2 U167 ( .A1(n146), .A2(n147), .ZN(\U7/Z_10 ) );
  NAND2_X2 U170 ( .A1(n148), .A2(n149), .ZN(\U7/Z_1 ) );
  NAND2_X2 U173 ( .A1(n150), .A2(n151), .ZN(\U7/Z_0 ) );
  NAND3_X2 U176 ( .A1(\add_46/A[0] ), .A2(n12), .A3(\add_46/A[1] ), .ZN(n40)
         );
  NOR4_X2 U181 ( .A1(n16), .A2(n13), .A3(\add_46/A[0] ), .A4(\add_46/A[2] ), 
        .ZN(n55) );
  OR3_X1 U196 ( .A1(FinalOutput[9]), .A2(FinalOutput[8]), .A3(FinalOutput[7]), 
        .ZN(n47) );
  OR3_X1 U197 ( .A1(FinalOutput[3]), .A2(FinalOutput[2]), .A3(FinalOutput[23]), 
        .ZN(n48) );
  OR3_X1 U198 ( .A1(FinalOutput[1]), .A2(FinalOutput[19]), .A3(FinalOutput[18]), .ZN(n49) );
  OR3_X1 U199 ( .A1(FinalOutput[14]), .A2(FinalOutput[13]), .A3(
        FinalOutput[12]), .ZN(n50) );
  OR3_X1 U200 ( .A1(\U13/DATA2_0 ), .A2(sig), .A3(n18), .ZN(n42) );
  DFF_X2 \addressI_reg[6]  ( .D(n396), .CK(clock), .Q(\add_54/A[6] ) );
  DFF_X2 \addressI_reg[5]  ( .D(n395), .CK(clock), .Q(\add_54/A[5] ) );
  DFF_X2 \addressI_reg[4]  ( .D(n394), .CK(clock), .Q(\add_54/A[4] ) );
  DFF_X2 \addressI_reg[3]  ( .D(n393), .CK(clock), .Q(\add_54/A[3] ) );
  DFF_X2 \addressI_reg[2]  ( .D(n392), .CK(clock), .Q(\add_54/A[2] ) );
  DFF_X2 \addressI_reg[1]  ( .D(n391), .CK(clock), .Q(\add_54/A[1] ) );
  DFF_X2 \addressI_reg[0]  ( .D(n153), .CK(clock), .Q(\add_54/A[0] ), .QN(n20)
         );
  DFF_X2 \addressI_reg[7]  ( .D(n152), .CK(clock), .Q(\add_54/A[7] ), .QN(n19)
         );
  AND4_X4 U3 ( .A1(n384), .A2(\add_46/A[0] ), .A3(n13), .A4(n12), .ZN(n386) );
  AND2_X4 U5 ( .A1(n23), .A2(n384), .ZN(n53) );
  NOR2_X4 U6 ( .A1(n16), .A2(n40), .ZN(n385) );
  INV_X4 U7 ( .A(n388), .ZN(n387) );
  AOI22_X2 U8 ( .A1(\U7/DATA3_0 ), .A2(n387), .B1(\U7/DATA2_0 ), .B2(n386), 
        .ZN(n150) );
  AOI22_X2 U9 ( .A1(\U7/DATA5_0 ), .A2(n53), .B1(\U7/DATA4_0 ), .B2(n385), 
        .ZN(n151) );
  AOI22_X2 U10 ( .A1(\U7/DATA3_1 ), .A2(n387), .B1(\U7/DATA2_1 ), .B2(n386), 
        .ZN(n148) );
  AOI22_X2 U11 ( .A1(\U7/DATA5_1 ), .A2(n53), .B1(\U7/DATA4_1 ), .B2(n385), 
        .ZN(n149) );
  AOI22_X2 U15 ( .A1(\U7/DATA3_2 ), .A2(n387), .B1(\U7/DATA2_2 ), .B2(n386), 
        .ZN(n126) );
  AOI22_X2 U16 ( .A1(\U7/DATA5_2 ), .A2(n53), .B1(\U7/DATA4_2 ), .B2(n385), 
        .ZN(n127) );
  AOI22_X2 U19 ( .A1(\U7/DATA3_3 ), .A2(n387), .B1(\U7/DATA2_3 ), .B2(n386), 
        .ZN(n104) );
  AOI22_X2 U20 ( .A1(\U7/DATA5_3 ), .A2(n53), .B1(\U7/DATA4_3 ), .B2(n385), 
        .ZN(n105) );
  AOI22_X2 U33 ( .A1(\U7/DATA3_4 ), .A2(n387), .B1(\U7/DATA2_4 ), .B2(n386), 
        .ZN(n81) );
  AOI22_X2 U34 ( .A1(\U7/DATA5_4 ), .A2(n53), .B1(\U7/DATA4_4 ), .B2(n385), 
        .ZN(n82) );
  AOI22_X2 U36 ( .A1(\U7/DATA3_5 ), .A2(n55), .B1(\U7/DATA2_5 ), .B2(n386), 
        .ZN(n63) );
  AOI22_X2 U37 ( .A1(\U7/DATA5_5 ), .A2(n53), .B1(\U7/DATA4_5 ), .B2(n385), 
        .ZN(n64) );
  AOI22_X2 U39 ( .A1(\U7/DATA3_6 ), .A2(n55), .B1(\U7/DATA2_6 ), .B2(n386), 
        .ZN(n61) );
  AOI22_X2 U40 ( .A1(\U7/DATA5_6 ), .A2(n53), .B1(\U7/DATA4_6 ), .B2(n385), 
        .ZN(n62) );
  AOI22_X2 U42 ( .A1(\U7/DATA3_7 ), .A2(n55), .B1(\U7/DATA2_7 ), .B2(n386), 
        .ZN(n59) );
  AOI22_X2 U43 ( .A1(\U7/DATA5_7 ), .A2(n53), .B1(\U7/DATA4_7 ), .B2(n385), 
        .ZN(n60) );
  AOI22_X2 U45 ( .A1(\U7/DATA3_8 ), .A2(n55), .B1(\U7/DATA2_8 ), .B2(n386), 
        .ZN(n57) );
  AOI22_X2 U46 ( .A1(\U7/DATA5_8 ), .A2(n53), .B1(\U7/DATA4_8 ), .B2(n385), 
        .ZN(n58) );
  AOI22_X2 U48 ( .A1(\U7/DATA3_9 ), .A2(n55), .B1(\U7/DATA2_9 ), .B2(n386), 
        .ZN(n51) );
  AOI22_X2 U49 ( .A1(\U7/DATA5_9 ), .A2(n53), .B1(\U7/DATA4_9 ), .B2(n385), 
        .ZN(n52) );
  AOI22_X2 U51 ( .A1(\U7/DATA3_10 ), .A2(n55), .B1(\U7/DATA2_10 ), .B2(n386), 
        .ZN(n146) );
  AOI22_X2 U52 ( .A1(\U7/DATA5_10 ), .A2(n53), .B1(\U7/DATA4_10 ), .B2(n385), 
        .ZN(n147) );
  AOI22_X2 U54 ( .A1(\U7/DATA3_11 ), .A2(n387), .B1(\U7/DATA2_11 ), .B2(n386), 
        .ZN(n144) );
  AOI22_X2 U55 ( .A1(\U7/DATA5_11 ), .A2(n53), .B1(\U7/DATA4_11 ), .B2(n385), 
        .ZN(n145) );
  AOI22_X2 U57 ( .A1(\U7/DATA3_12 ), .A2(n387), .B1(\U7/DATA2_12 ), .B2(n386), 
        .ZN(n142) );
  AOI22_X2 U58 ( .A1(\U7/DATA5_12 ), .A2(n53), .B1(\U7/DATA4_12 ), .B2(n385), 
        .ZN(n143) );
  AOI22_X2 U60 ( .A1(\U7/DATA3_13 ), .A2(n55), .B1(\U7/DATA2_13 ), .B2(n386), 
        .ZN(n140) );
  AOI22_X2 U61 ( .A1(\U7/DATA5_13 ), .A2(n53), .B1(\U7/DATA4_13 ), .B2(n385), 
        .ZN(n141) );
  AOI22_X2 U63 ( .A1(\U7/DATA3_14 ), .A2(n387), .B1(\U7/DATA2_14 ), .B2(n386), 
        .ZN(n138) );
  AOI22_X2 U64 ( .A1(\U7/DATA5_14 ), .A2(n53), .B1(\U7/DATA4_14 ), .B2(n385), 
        .ZN(n139) );
  AOI22_X2 U66 ( .A1(\U7/DATA3_15 ), .A2(n387), .B1(\U7/DATA2_15 ), .B2(n386), 
        .ZN(n136) );
  AOI22_X2 U67 ( .A1(\U7/DATA5_15 ), .A2(n53), .B1(\U7/DATA4_15 ), .B2(n385), 
        .ZN(n137) );
  AOI22_X2 U69 ( .A1(\U7/DATA3_16 ), .A2(n55), .B1(\U7/DATA2_16 ), .B2(n386), 
        .ZN(n134) );
  AOI22_X2 U70 ( .A1(\U7/DATA5_16 ), .A2(n53), .B1(\U7/DATA4_16 ), .B2(n385), 
        .ZN(n135) );
  AOI22_X2 U72 ( .A1(\U7/DATA3_17 ), .A2(n55), .B1(\U7/DATA2_17 ), .B2(n386), 
        .ZN(n132) );
  AOI22_X2 U73 ( .A1(\U7/DATA5_17 ), .A2(n53), .B1(\U7/DATA4_17 ), .B2(n385), 
        .ZN(n133) );
  AOI22_X2 U75 ( .A1(\U7/DATA3_18 ), .A2(n55), .B1(\U7/DATA2_18 ), .B2(n386), 
        .ZN(n130) );
  AOI22_X2 U76 ( .A1(\U7/DATA5_18 ), .A2(n53), .B1(\U7/DATA4_18 ), .B2(n385), 
        .ZN(n131) );
  AOI22_X2 U78 ( .A1(\U7/DATA3_19 ), .A2(n55), .B1(\U7/DATA2_19 ), .B2(n386), 
        .ZN(n128) );
  AOI22_X2 U79 ( .A1(\U7/DATA5_19 ), .A2(n53), .B1(\U7/DATA4_19 ), .B2(n385), 
        .ZN(n129) );
  AOI22_X2 U81 ( .A1(\U7/DATA3_20 ), .A2(n387), .B1(\U7/DATA2_20 ), .B2(n386), 
        .ZN(n124) );
  AOI22_X2 U82 ( .A1(\U7/DATA5_20 ), .A2(n53), .B1(\U7/DATA4_20 ), .B2(n385), 
        .ZN(n125) );
  AOI22_X2 U84 ( .A1(\U7/DATA3_21 ), .A2(n387), .B1(\U7/DATA2_21 ), .B2(n386), 
        .ZN(n122) );
  AOI22_X2 U85 ( .A1(\U7/DATA5_21 ), .A2(n53), .B1(\U7/DATA4_21 ), .B2(n385), 
        .ZN(n123) );
  AOI22_X2 U87 ( .A1(\U7/DATA3_22 ), .A2(n387), .B1(\U7/DATA2_22 ), .B2(n386), 
        .ZN(n120) );
  AOI22_X2 U88 ( .A1(\U7/DATA5_22 ), .A2(n53), .B1(\U7/DATA4_22 ), .B2(n385), 
        .ZN(n121) );
  AOI22_X2 U90 ( .A1(\U7/DATA3_23 ), .A2(n387), .B1(\U7/DATA2_23 ), .B2(n386), 
        .ZN(n118) );
  AOI22_X2 U91 ( .A1(\U7/DATA5_23 ), .A2(n53), .B1(\U7/DATA4_23 ), .B2(n385), 
        .ZN(n119) );
  AOI22_X2 U93 ( .A1(\U7/DATA3_24 ), .A2(n387), .B1(\U7/DATA2_24 ), .B2(n386), 
        .ZN(n116) );
  AOI22_X2 U94 ( .A1(\U7/DATA5_24 ), .A2(n53), .B1(\U7/DATA4_24 ), .B2(n385), 
        .ZN(n117) );
  AOI22_X2 U96 ( .A1(\U7/DATA3_25 ), .A2(n387), .B1(\U7/DATA2_25 ), .B2(n386), 
        .ZN(n114) );
  AOI22_X2 U97 ( .A1(\U7/DATA5_25 ), .A2(n53), .B1(\U7/DATA4_25 ), .B2(n385), 
        .ZN(n115) );
  AOI22_X2 U99 ( .A1(\U7/DATA3_26 ), .A2(n387), .B1(\U7/DATA2_26 ), .B2(n386), 
        .ZN(n112) );
  AOI22_X2 U100 ( .A1(\U7/DATA5_26 ), .A2(n53), .B1(\U7/DATA4_26 ), .B2(n385), 
        .ZN(n113) );
  AOI22_X2 U102 ( .A1(\U7/DATA3_27 ), .A2(n387), .B1(\U7/DATA2_27 ), .B2(n386), 
        .ZN(n110) );
  AOI22_X2 U103 ( .A1(\U7/DATA5_27 ), .A2(n53), .B1(\U7/DATA4_27 ), .B2(n385), 
        .ZN(n111) );
  AOI22_X2 U105 ( .A1(\U7/DATA3_28 ), .A2(n387), .B1(\U7/DATA2_28 ), .B2(n386), 
        .ZN(n108) );
  AOI22_X2 U106 ( .A1(\U7/DATA5_28 ), .A2(n53), .B1(\U7/DATA4_28 ), .B2(n385), 
        .ZN(n109) );
  AOI22_X2 U108 ( .A1(\U7/DATA3_29 ), .A2(n387), .B1(\U7/DATA2_29 ), .B2(n386), 
        .ZN(n106) );
  AOI22_X2 U109 ( .A1(\U7/DATA5_29 ), .A2(n53), .B1(\U7/DATA4_29 ), .B2(n385), 
        .ZN(n107) );
  AOI22_X2 U111 ( .A1(\U7/DATA3_30 ), .A2(n387), .B1(\U7/DATA2_30 ), .B2(n386), 
        .ZN(n102) );
  AOI22_X2 U112 ( .A1(\U7/DATA5_30 ), .A2(n53), .B1(\U7/DATA4_30 ), .B2(n385), 
        .ZN(n103) );
  AOI22_X2 U114 ( .A1(\U7/DATA3_31 ), .A2(n387), .B1(\U7/DATA2_31 ), .B2(n386), 
        .ZN(n100) );
  AOI22_X2 U115 ( .A1(\U7/DATA5_31 ), .A2(n53), .B1(\U7/DATA4_31 ), .B2(n385), 
        .ZN(n101) );
  AOI22_X2 U117 ( .A1(\U7/DATA3_32 ), .A2(n387), .B1(\U7/DATA2_32 ), .B2(n386), 
        .ZN(n98) );
  AOI22_X2 U118 ( .A1(\U7/DATA5_32 ), .A2(n53), .B1(\U7/DATA4_32 ), .B2(n385), 
        .ZN(n99) );
  AOI22_X2 U120 ( .A1(\U7/DATA3_33 ), .A2(n387), .B1(\U7/DATA2_33 ), .B2(n386), 
        .ZN(n95) );
  AOI22_X2 U121 ( .A1(\U7/DATA5_33 ), .A2(n53), .B1(\U7/DATA4_33 ), .B2(n385), 
        .ZN(n97) );
  AOI22_X2 U123 ( .A1(\U7/DATA3_34 ), .A2(n55), .B1(\U7/DATA2_34 ), .B2(n386), 
        .ZN(n93) );
  AOI22_X2 U124 ( .A1(\U7/DATA5_34 ), .A2(n53), .B1(\U7/DATA4_34 ), .B2(n385), 
        .ZN(n94) );
  AOI22_X2 U126 ( .A1(\U7/DATA3_35 ), .A2(n55), .B1(\U7/DATA2_35 ), .B2(n386), 
        .ZN(n91) );
  AOI22_X2 U127 ( .A1(\U7/DATA5_35 ), .A2(n53), .B1(\U7/DATA4_35 ), .B2(n385), 
        .ZN(n92) );
  AOI22_X2 U129 ( .A1(\U7/DATA3_36 ), .A2(n55), .B1(\U7/DATA2_36 ), .B2(n386), 
        .ZN(n89) );
  AOI22_X2 U130 ( .A1(\U7/DATA5_36 ), .A2(n53), .B1(\U7/DATA4_36 ), .B2(n385), 
        .ZN(n90) );
  AOI22_X2 U132 ( .A1(\U7/DATA3_37 ), .A2(n55), .B1(\U7/DATA2_37 ), .B2(n386), 
        .ZN(n87) );
  AOI22_X2 U133 ( .A1(\U7/DATA5_37 ), .A2(n53), .B1(\U7/DATA4_37 ), .B2(n385), 
        .ZN(n88) );
  AOI22_X2 U135 ( .A1(\U7/DATA3_38 ), .A2(n55), .B1(\U7/DATA2_38 ), .B2(n386), 
        .ZN(n85) );
  AOI22_X2 U136 ( .A1(\U7/DATA5_38 ), .A2(n53), .B1(\U7/DATA4_38 ), .B2(n385), 
        .ZN(n86) );
  AOI22_X2 U138 ( .A1(\U7/DATA3_39 ), .A2(n55), .B1(\U7/DATA2_39 ), .B2(n386), 
        .ZN(n83) );
  AOI22_X2 U139 ( .A1(\U7/DATA5_39 ), .A2(n53), .B1(\U7/DATA4_39 ), .B2(n385), 
        .ZN(n84) );
  AOI22_X2 U141 ( .A1(\U7/DATA3_40 ), .A2(n55), .B1(\U7/DATA2_40 ), .B2(n386), 
        .ZN(n79) );
  AOI22_X2 U142 ( .A1(\U7/DATA5_40 ), .A2(n53), .B1(\U7/DATA4_40 ), .B2(n385), 
        .ZN(n80) );
  AOI22_X2 U144 ( .A1(\U7/DATA3_41 ), .A2(n55), .B1(\U7/DATA2_41 ), .B2(n386), 
        .ZN(n77) );
  AOI22_X2 U145 ( .A1(\U7/DATA5_41 ), .A2(n53), .B1(\U7/DATA4_41 ), .B2(n385), 
        .ZN(n78) );
  AOI22_X2 U147 ( .A1(\U7/DATA3_42 ), .A2(n55), .B1(\U7/DATA2_42 ), .B2(n386), 
        .ZN(n75) );
  AOI22_X2 U148 ( .A1(\U7/DATA5_42 ), .A2(n53), .B1(\U7/DATA4_42 ), .B2(n385), 
        .ZN(n76) );
  AOI22_X2 U150 ( .A1(\U7/DATA3_43 ), .A2(n387), .B1(\U7/DATA2_43 ), .B2(n386), 
        .ZN(n73) );
  AOI22_X2 U151 ( .A1(\U7/DATA5_43 ), .A2(n53), .B1(\U7/DATA4_43 ), .B2(n385), 
        .ZN(n74) );
  AOI22_X2 U153 ( .A1(\U7/DATA3_44 ), .A2(n387), .B1(\U7/DATA2_44 ), .B2(n386), 
        .ZN(n71) );
  AOI22_X2 U154 ( .A1(\U7/DATA5_44 ), .A2(n53), .B1(\U7/DATA4_44 ), .B2(n385), 
        .ZN(n72) );
  AOI22_X2 U156 ( .A1(\U7/DATA3_45 ), .A2(n387), .B1(\U7/DATA2_45 ), .B2(n386), 
        .ZN(n69) );
  AOI22_X2 U157 ( .A1(\U7/DATA5_45 ), .A2(n53), .B1(\U7/DATA4_45 ), .B2(n385), 
        .ZN(n70) );
  AOI22_X2 U159 ( .A1(\U7/DATA3_46 ), .A2(n387), .B1(\U7/DATA2_46 ), .B2(n386), 
        .ZN(n67) );
  AOI22_X2 U160 ( .A1(\U7/DATA5_46 ), .A2(n53), .B1(\U7/DATA4_46 ), .B2(n385), 
        .ZN(n68) );
  AOI22_X2 U162 ( .A1(\U7/DATA3_47 ), .A2(n387), .B1(\U7/DATA2_47 ), .B2(n386), 
        .ZN(n65) );
  AOI22_X2 U163 ( .A1(\U7/DATA5_47 ), .A2(n53), .B1(\U7/DATA4_47 ), .B2(n385), 
        .ZN(n66) );
  AOI21_X2 U165 ( .B1(n37), .B2(n13), .A(n38), .ZN(n39) );
  AOI22_X1 U166 ( .A1(\U4/DATA1_6 ), .A2(n23), .B1(\add_54/A[6] ), .B2(n26), 
        .ZN(n25) );
  AOI22_X1 U168 ( .A1(\U4/DATA1_4 ), .A2(n23), .B1(\add_54/A[4] ), .B2(n26), 
        .ZN(n28) );
  AOI22_X1 U169 ( .A1(\U4/DATA1_3 ), .A2(n23), .B1(\add_54/A[3] ), .B2(n26), 
        .ZN(n29) );
  AOI22_X1 U171 ( .A1(\U4/DATA1_2 ), .A2(n23), .B1(\add_54/A[2] ), .B2(n26), 
        .ZN(n30) );
  AOI22_X1 U172 ( .A1(\U4/DATA1_1 ), .A2(n23), .B1(\add_54/A[1] ), .B2(n26), 
        .ZN(n31) );
  OAI21_X2 U174 ( .B1(\add_46/A[0] ), .B2(n400), .A(n32), .ZN(n38) );
  AOI22_X1 U175 ( .A1(\U4/DATA1_5 ), .A2(n23), .B1(\add_54/A[5] ), .B2(n26), 
        .ZN(n27) );
  INV_X4 U177 ( .A(n55), .ZN(n388) );
  NOR3_X2 U178 ( .A1(\add_46/A[0] ), .A2(\add_46/A[1] ), .A3(n12), .ZN(n23) );
  OAI21_X2 U179 ( .B1(n389), .B2(n19), .A(n22), .ZN(n152) );
  OAI21_X2 U180 ( .B1(n401), .B2(\add_54/carry[7] ), .A(n390), .ZN(n24) );
  OAI21_X2 U182 ( .B1(n34), .B2(\add_46/A[0] ), .A(n35), .ZN(n33) );
  OAI21_X2 U183 ( .B1(n397), .B2(n13), .A(n36), .ZN(n155) );
  INV_X4 U184 ( .A(n24), .ZN(n389) );
  INV_X4 U185 ( .A(n26), .ZN(n390) );
  INV_X4 U186 ( .A(n31), .ZN(n391) );
  INV_X4 U187 ( .A(n30), .ZN(n392) );
  INV_X4 U188 ( .A(n29), .ZN(n393) );
  INV_X4 U189 ( .A(n28), .ZN(n394) );
  INV_X4 U190 ( .A(n27), .ZN(n395) );
  INV_X4 U191 ( .A(n25), .ZN(n396) );
  INV_X4 U192 ( .A(n38), .ZN(n397) );
  INV_X4 U193 ( .A(n35), .ZN(n398) );
  INV_X4 U194 ( .A(n33), .ZN(n399) );
  INV_X4 U195 ( .A(n37), .ZN(n400) );
  INV_X4 U201 ( .A(n23), .ZN(n401) );
  INV_X4 U202 ( .A(sig), .ZN(n402) );
endmodule


module write_enable ( input_data, input_data2, signal, signal2 );
  input [47:0] input_data;
  input [47:0] input_data2;
  output signal, signal2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  NAND4_X2 U1 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(n4) );
  NAND4_X2 U6 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n3) );
  NAND4_X2 U11 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(n2) );
  NAND4_X2 U16 ( .A1(n17), .A2(n18), .A3(n19), .A4(n20), .ZN(n1) );
  NAND4_X2 U21 ( .A1(n25), .A2(n26), .A3(n27), .A4(n28), .ZN(n24) );
  NOR3_X2 U22 ( .A1(input_data[39]), .A2(input_data[40]), .A3(input_data[3]), 
        .ZN(n28) );
  NOR3_X2 U23 ( .A1(input_data[36]), .A2(input_data[38]), .A3(input_data[37]), 
        .ZN(n27) );
  NOR3_X2 U24 ( .A1(input_data[33]), .A2(input_data[35]), .A3(input_data[34]), 
        .ZN(n26) );
  NOR3_X2 U25 ( .A1(input_data[30]), .A2(input_data[32]), .A3(input_data[31]), 
        .ZN(n25) );
  NAND4_X2 U26 ( .A1(n29), .A2(n30), .A3(n31), .A4(n32), .ZN(n23) );
  NOR3_X2 U27 ( .A1(input_data[7]), .A2(input_data[9]), .A3(input_data[8]), 
        .ZN(n32) );
  NOR3_X2 U28 ( .A1(input_data[4]), .A2(input_data[6]), .A3(input_data[5]), 
        .ZN(n31) );
  NOR3_X2 U29 ( .A1(input_data[44]), .A2(input_data[46]), .A3(input_data[45]), 
        .ZN(n30) );
  NOR3_X2 U30 ( .A1(input_data[41]), .A2(input_data[43]), .A3(input_data[42]), 
        .ZN(n29) );
  NAND4_X2 U31 ( .A1(n33), .A2(n34), .A3(n35), .A4(n36), .ZN(n22) );
  NOR3_X2 U32 ( .A1(input_data[17]), .A2(input_data[19]), .A3(input_data[18]), 
        .ZN(n36) );
  NOR3_X2 U33 ( .A1(input_data[14]), .A2(input_data[16]), .A3(input_data[15]), 
        .ZN(n35) );
  NOR3_X2 U34 ( .A1(input_data[11]), .A2(input_data[13]), .A3(input_data[12]), 
        .ZN(n34) );
  NOR2_X2 U35 ( .A1(input_data[10]), .A2(input_data[0]), .ZN(n33) );
  NAND4_X2 U36 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(n21) );
  NOR3_X2 U37 ( .A1(input_data[28]), .A2(input_data[2]), .A3(input_data[29]), 
        .ZN(n40) );
  NOR3_X2 U38 ( .A1(input_data[25]), .A2(input_data[27]), .A3(input_data[26]), 
        .ZN(n39) );
  NOR3_X2 U39 ( .A1(input_data[22]), .A2(input_data[24]), .A3(input_data[23]), 
        .ZN(n38) );
  NOR3_X2 U40 ( .A1(input_data[1]), .A2(input_data[21]), .A3(input_data[20]), 
        .ZN(n37) );
  OR4_X1 U41 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(signal2) );
  OR4_X1 U42 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(signal) );
  NOR2_X1 U2 ( .A1(input_data2[10]), .A2(input_data2[0]), .ZN(n13) );
  NOR3_X1 U3 ( .A1(input_data2[41]), .A2(input_data2[43]), .A3(input_data2[42]), .ZN(n9) );
  NOR3_X1 U4 ( .A1(input_data2[30]), .A2(input_data2[32]), .A3(input_data2[31]), .ZN(n5) );
  NOR3_X1 U5 ( .A1(input_data2[11]), .A2(input_data2[13]), .A3(input_data2[12]), .ZN(n14) );
  NOR3_X1 U7 ( .A1(input_data2[1]), .A2(input_data2[21]), .A3(input_data2[20]), 
        .ZN(n17) );
  NOR3_X1 U8 ( .A1(input_data2[44]), .A2(input_data2[46]), .A3(input_data2[45]), .ZN(n10) );
  NOR3_X1 U9 ( .A1(input_data2[39]), .A2(input_data2[40]), .A3(input_data2[3]), 
        .ZN(n8) );
  NOR3_X1 U10 ( .A1(input_data2[36]), .A2(input_data2[38]), .A3(
        input_data2[37]), .ZN(n7) );
  NOR3_X1 U12 ( .A1(input_data2[33]), .A2(input_data2[35]), .A3(
        input_data2[34]), .ZN(n6) );
  NOR3_X1 U13 ( .A1(input_data2[28]), .A2(input_data2[2]), .A3(input_data2[29]), .ZN(n20) );
  NOR3_X1 U14 ( .A1(input_data2[25]), .A2(input_data2[27]), .A3(
        input_data2[26]), .ZN(n19) );
  NOR3_X1 U15 ( .A1(input_data2[22]), .A2(input_data2[24]), .A3(
        input_data2[23]), .ZN(n18) );
  NOR3_X1 U17 ( .A1(input_data2[7]), .A2(input_data2[9]), .A3(input_data2[8]), 
        .ZN(n12) );
  NOR3_X1 U18 ( .A1(input_data2[4]), .A2(input_data2[6]), .A3(input_data2[5]), 
        .ZN(n11) );
  NOR3_X1 U19 ( .A1(input_data2[17]), .A2(input_data2[19]), .A3(
        input_data2[18]), .ZN(n16) );
  NOR3_X1 U20 ( .A1(input_data2[14]), .A2(input_data2[16]), .A3(
        input_data2[15]), .ZN(n15) );
endmodule


module v_sched ( signal, signal2, clock, reset, write_addr1, we1, write_addr2, 
        we2, write_addr3, we3, write_addr4, we4, sig_I, count2 );
  output [8:0] write_addr1;
  output [8:0] write_addr2;
  output [8:0] write_addr3;
  output [8:0] write_addr4;
  input signal, signal2, clock, reset, sig_I, count2;
  output we1, we2, we3, we4;
  wire   \U20/DATA2_0 , \U6/DATA1_1 , \U6/DATA1_2 , \U6/DATA1_3 , \U6/DATA1_4 ,
         \U6/DATA1_5 , \U6/DATA1_6 , \U6/DATA1_7 , \mult_add_42_aco/a[2] ,
         \mult_add_42_aco/a[1] , \mult_add_42_aco/a[0] , \r344/carry[8] ,
         \r344/carry[7] , \r344/carry[6] , \r344/carry[5] , \r344/carry[4] ,
         \r344/carry[3] , \r344/carry[2] , n16, n17, n18, n19, n20, n21, n22,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n193, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235;
  assign \U20/DATA2_0  = reset;

  HA_X1 \r344/U1_1_1  ( .A(write_addr3[1]), .B(write_addr3[0]), .CO(
        \r344/carry[2] ), .S(\U6/DATA1_1 ) );
  HA_X1 \r344/U1_1_2  ( .A(write_addr3[2]), .B(\r344/carry[2] ), .CO(
        \r344/carry[3] ), .S(\U6/DATA1_2 ) );
  HA_X1 \r344/U1_1_3  ( .A(write_addr3[3]), .B(\r344/carry[3] ), .CO(
        \r344/carry[4] ), .S(\U6/DATA1_3 ) );
  HA_X1 \r344/U1_1_4  ( .A(write_addr3[4]), .B(\r344/carry[4] ), .CO(
        \r344/carry[5] ), .S(\U6/DATA1_4 ) );
  HA_X1 \r344/U1_1_5  ( .A(write_addr3[5]), .B(\r344/carry[5] ), .CO(
        \r344/carry[6] ), .S(\U6/DATA1_5 ) );
  HA_X1 \r344/U1_1_6  ( .A(write_addr3[6]), .B(\r344/carry[6] ), .CO(
        \r344/carry[7] ), .S(\U6/DATA1_6 ) );
  HA_X1 \r344/U1_1_7  ( .A(write_addr3[7]), .B(\r344/carry[7] ), .CO(
        \r344/carry[8] ), .S(\U6/DATA1_7 ) );
  DFF_X1 \count_reg[0]  ( .D(n63), .CK(clock), .Q(\mult_add_42_aco/a[0] ), 
        .QN(n18) );
  DFF_X1 \count_reg[2]  ( .D(n62), .CK(clock), .Q(\mult_add_42_aco/a[2] ), 
        .QN(n16) );
  DFF_X1 \count_reg[1]  ( .D(n61), .CK(clock), .Q(\mult_add_42_aco/a[1] ), 
        .QN(n17) );
  OAI221_X2 U11 ( .B1(n36), .B2(n37), .C1(count2), .C2(n235), .A(n38), .ZN(n34) );
  NAND3_X2 U12 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n38) );
  NOR2_X2 U13 ( .A1(n234), .A2(n40), .ZN(n36) );
  XOR2_X2 U14 ( .A(write_addr3[8]), .B(\r344/carry[8] ), .Z(n40) );
  OAI22_X2 U18 ( .A1(n43), .A2(n21), .B1(n230), .B2(n44), .ZN(n57) );
  OAI22_X2 U20 ( .A1(n45), .A2(n20), .B1(n231), .B2(n46), .ZN(n58) );
  OAI22_X2 U22 ( .A1(n47), .A2(n19), .B1(n232), .B2(n48), .ZN(n59) );
  NAND4_X2 U25 ( .A1(n51), .A2(n46), .A3(n48), .A4(n44), .ZN(n50) );
  NAND3_X2 U26 ( .A1(\mult_add_42_aco/a[1] ), .A2(n16), .A3(
        \mult_add_42_aco/a[0] ), .ZN(n44) );
  NAND3_X2 U27 ( .A1(n18), .A2(n16), .A3(\mult_add_42_aco/a[1] ), .ZN(n46) );
  NAND3_X2 U30 ( .A1(n17), .A2(n16), .A3(\mult_add_42_aco/a[0] ), .ZN(n48) );
  NAND2_X2 U31 ( .A1(n52), .A2(n235), .ZN(n37) );
  NAND3_X2 U33 ( .A1(\mult_add_42_aco/a[0] ), .A2(n17), .A3(n41), .ZN(n54) );
  NAND3_X2 U34 ( .A1(\mult_add_42_aco/a[1] ), .A2(n18), .A3(n41), .ZN(n53) );
  NAND3_X2 U36 ( .A1(\mult_add_42_aco/a[0] ), .A2(\mult_add_42_aco/a[1] ), 
        .A3(n41), .ZN(n55) );
  OAI22_X2 U37 ( .A1(n18), .A2(n35), .B1(\mult_add_42_aco/a[0] ), .B2(n233), 
        .ZN(n63) );
  NOR2_X2 U38 ( .A1(n56), .A2(\mult_add_42_aco/a[0] ), .ZN(n39) );
  NOR2_X2 U39 ( .A1(n52), .A2(sig_I), .ZN(n41) );
  OAI221_X2 U40 ( .B1(n16), .B2(n17), .C1(n56), .C2(n18), .A(signal), .ZN(n52)
         );
  NAND2_X2 U41 ( .A1(\mult_add_42_aco/a[2] ), .A2(n17), .ZN(n56) );
  OR4_X1 U58 ( .A1(n41), .A2(n39), .A3(sig_I), .A4(\U20/DATA2_0 ), .ZN(n35) );
  DFF_X2 \addressV_reg[1]  ( .D(n222), .CK(clock), .Q(write_addr3[1]) );
  DFF_X2 \addressV_reg[2]  ( .D(n223), .CK(clock), .Q(write_addr3[2]) );
  DFF_X2 \addressV_reg[3]  ( .D(n224), .CK(clock), .Q(write_addr3[3]) );
  DFF_X2 \addressV_reg[4]  ( .D(n225), .CK(clock), .Q(write_addr3[4]) );
  DFF_X2 \addressV_reg[5]  ( .D(n226), .CK(clock), .Q(write_addr3[5]) );
  DFF_X2 \addressV_reg[6]  ( .D(n227), .CK(clock), .Q(write_addr3[6]) );
  DFF_X2 \addressV_reg[7]  ( .D(n228), .CK(clock), .Q(write_addr3[7]) );
  DFF_X2 \addressV_reg[8]  ( .D(n229), .CK(clock), .Q(write_addr3[8]) );
  DFF_X2 we1_reg ( .D(n60), .CK(clock), .Q(we1), .QN(n193) );
  DFF_X2 we3_reg ( .D(n58), .CK(clock), .Q(we3), .QN(n20) );
  DFF_X2 we2_reg ( .D(n59), .CK(clock), .Q(we2), .QN(n19) );
  DFF_X2 we4_reg ( .D(n57), .CK(clock), .Q(we4), .QN(n21) );
  DFF_X2 \addressV_reg[0]  ( .D(n221), .CK(clock), .Q(write_addr3[0]), .QN(n22) );
  OAI21_X2 U3 ( .B1(n193), .B2(n51), .A(n50), .ZN(n60) );
  AOI21_X2 U4 ( .B1(n233), .B2(n37), .A(n234), .ZN(n25) );
  OAI21_X2 U5 ( .B1(n39), .B2(n233), .A(n35), .ZN(n26) );
  OAI21_X2 U6 ( .B1(n37), .B2(n48), .A(n233), .ZN(n51) );
  AOI22_X2 U7 ( .A1(n34), .A2(n35), .B1(write_addr3[8]), .B2(n26), .ZN(n33) );
  OAI21_X2 U8 ( .B1(n37), .B2(n44), .A(n233), .ZN(n45) );
  OAI21_X2 U9 ( .B1(n37), .B2(n46), .A(n233), .ZN(n47) );
  OAI211_X2 U10 ( .C1(n17), .C2(n35), .A(n53), .B(n54), .ZN(n61) );
  OAI21_X2 U15 ( .B1(n16), .B2(n35), .A(n55), .ZN(n62) );
  AOI22_X2 U16 ( .A1(\U6/DATA1_7 ), .A2(n25), .B1(write_addr3[7]), .B2(n26), 
        .ZN(n24) );
  AOI22_X2 U17 ( .A1(\U6/DATA1_6 ), .A2(n25), .B1(write_addr3[6]), .B2(n26), 
        .ZN(n27) );
  AOI22_X2 U19 ( .A1(\U6/DATA1_5 ), .A2(n25), .B1(write_addr3[5]), .B2(n26), 
        .ZN(n28) );
  AOI22_X2 U21 ( .A1(\U6/DATA1_4 ), .A2(n25), .B1(write_addr3[4]), .B2(n26), 
        .ZN(n29) );
  AOI22_X2 U23 ( .A1(\U6/DATA1_3 ), .A2(n25), .B1(write_addr3[3]), .B2(n26), 
        .ZN(n30) );
  AOI22_X2 U24 ( .A1(\U6/DATA1_2 ), .A2(n25), .B1(write_addr3[2]), .B2(n26), 
        .ZN(n31) );
  AOI22_X2 U28 ( .A1(\U6/DATA1_1 ), .A2(n25), .B1(write_addr3[1]), .B2(n26), 
        .ZN(n32) );
  AOI22_X2 U29 ( .A1(n26), .A2(write_addr3[0]), .B1(n22), .B2(n25), .ZN(n42)
         );
  OAI21_X2 U32 ( .B1(n234), .B2(n37), .A(n233), .ZN(n43) );
  BUF_X4 U35 ( .A(write_addr3[8]), .Z(write_addr2[8]) );
  BUF_X4 U42 ( .A(write_addr3[8]), .Z(write_addr1[8]) );
  BUF_X4 U43 ( .A(write_addr3[8]), .Z(write_addr4[8]) );
  BUF_X4 U44 ( .A(write_addr3[7]), .Z(write_addr2[7]) );
  BUF_X4 U45 ( .A(write_addr3[7]), .Z(write_addr1[7]) );
  BUF_X4 U46 ( .A(write_addr3[7]), .Z(write_addr4[7]) );
  BUF_X4 U47 ( .A(write_addr3[6]), .Z(write_addr2[6]) );
  BUF_X4 U48 ( .A(write_addr3[6]), .Z(write_addr1[6]) );
  BUF_X4 U49 ( .A(write_addr3[6]), .Z(write_addr4[6]) );
  BUF_X4 U50 ( .A(write_addr3[5]), .Z(write_addr2[5]) );
  BUF_X4 U51 ( .A(write_addr3[5]), .Z(write_addr1[5]) );
  BUF_X4 U52 ( .A(write_addr3[5]), .Z(write_addr4[5]) );
  BUF_X4 U53 ( .A(write_addr3[4]), .Z(write_addr2[4]) );
  BUF_X4 U54 ( .A(write_addr3[4]), .Z(write_addr1[4]) );
  BUF_X4 U55 ( .A(write_addr3[4]), .Z(write_addr4[4]) );
  BUF_X4 U56 ( .A(write_addr3[3]), .Z(write_addr2[3]) );
  BUF_X4 U57 ( .A(write_addr3[3]), .Z(write_addr1[3]) );
  BUF_X4 U59 ( .A(write_addr3[3]), .Z(write_addr4[3]) );
  BUF_X4 U60 ( .A(write_addr3[2]), .Z(write_addr2[2]) );
  BUF_X4 U61 ( .A(write_addr3[2]), .Z(write_addr1[2]) );
  BUF_X4 U62 ( .A(write_addr3[2]), .Z(write_addr4[2]) );
  BUF_X4 U63 ( .A(write_addr3[1]), .Z(write_addr2[1]) );
  BUF_X4 U64 ( .A(write_addr3[1]), .Z(write_addr1[1]) );
  BUF_X4 U65 ( .A(write_addr3[1]), .Z(write_addr4[1]) );
  BUF_X4 U66 ( .A(write_addr3[0]), .Z(write_addr2[0]) );
  BUF_X4 U67 ( .A(write_addr3[0]), .Z(write_addr1[0]) );
  BUF_X4 U68 ( .A(write_addr3[0]), .Z(write_addr4[0]) );
  INV_X4 U69 ( .A(n42), .ZN(n221) );
  INV_X4 U70 ( .A(n32), .ZN(n222) );
  INV_X4 U71 ( .A(n31), .ZN(n223) );
  INV_X4 U72 ( .A(n30), .ZN(n224) );
  INV_X4 U73 ( .A(n29), .ZN(n225) );
  INV_X4 U74 ( .A(n28), .ZN(n226) );
  INV_X4 U75 ( .A(n27), .ZN(n227) );
  INV_X4 U76 ( .A(n24), .ZN(n228) );
  INV_X4 U77 ( .A(n33), .ZN(n229) );
  INV_X4 U78 ( .A(n43), .ZN(n230) );
  INV_X4 U79 ( .A(n45), .ZN(n231) );
  INV_X4 U80 ( .A(n47), .ZN(n232) );
  INV_X4 U81 ( .A(n41), .ZN(n233) );
  INV_X4 U82 ( .A(n39), .ZN(n234) );
  INV_X4 U83 ( .A(sig_I), .ZN(n235) );
endmodule


module top_4 ( clock, reset, Vout, mult_output, vop1, vop2, vop3, vop4, 
        Rowread1, Rowread2, Rowread3, Rowread4, we1, we2, we3, we4, 
        write_addr1, write_addr2, write_addr3, write_addr4, op_reg, outI, 
        addressI, SyncMultY, SyncV, op1, subOut, multinput, op_final, dataI, 
        delay1, adder_out7, adder_out7_imag, adder_out1, adder_out2, 
        adder_out1_imag, adder_out2_imag, accum_output, accum_input, 
        adder_input, accum_output_imag, accum_input_imag, adder_input_imag, 
        div_output, diagonalC, diagonalD, adder_out3, adder_out4, 
        adder_out3_imag, adder_out4_imag, X, Y, EnableChange, NewElement, 
        ReadAddress1, ReadAddress2, WE, WriteReq, WriteBus, ReadBus1, ReadBus2, 
        SubOutput, AddOutput, AddInput1, AddInput2, SubInput1, SubInput2, 
        EOC_Flag, sig_OP, diagOut, Mul_In );
  output [47:0] Vout;
  output [48:0] mult_output;
  input [47:0] vop1;
  input [47:0] vop2;
  input [47:0] vop3;
  input [47:0] vop4;
  output [8:0] Rowread1;
  output [8:0] Rowread2;
  output [8:0] Rowread3;
  output [8:0] Rowread4;
  output [8:0] write_addr1;
  output [8:0] write_addr2;
  output [8:0] write_addr3;
  output [8:0] write_addr4;
  output [47:0] op_reg;
  input [191:0] outI;
  output [7:0] addressI;
  output [47:0] SyncMultY;
  output [47:0] SyncV;
  output [47:0] op1;
  input [47:0] subOut;
  input [47:0] multinput;
  input [47:0] op_final;
  output [47:0] dataI;
  output [47:0] delay1;
  input [23:0] adder_out7;
  input [23:0] adder_out7_imag;
  output [23:0] adder_out1;
  output [23:0] adder_out2;
  output [23:0] adder_out1_imag;
  output [23:0] adder_out2_imag;
  input [23:0] accum_output;
  output [23:0] accum_input;
  output [23:0] adder_input;
  input [23:0] accum_output_imag;
  output [23:0] accum_input_imag;
  output [23:0] adder_input_imag;
  input [47:0] div_output;
  output [23:0] diagonalC;
  output [23:0] diagonalD;
  output [23:0] adder_out3;
  output [23:0] adder_out4;
  output [23:0] adder_out3_imag;
  output [23:0] adder_out4_imag;
  input [15:0] X;
  input [15:0] Y;
  input [47:0] NewElement;
  output [10:0] ReadAddress1;
  output [10:0] ReadAddress2;
  output [10:0] WriteReq;
  output [255:0] WriteBus;
  input [255:0] ReadBus1;
  input [255:0] ReadBus2;
  input [23:0] SubOutput;
  input [23:0] AddOutput;
  output [23:0] AddInput1;
  output [23:0] AddInput2;
  output [23:0] SubInput1;
  output [23:0] SubInput2;
  output [47:0] diagOut;
  output [47:0] Mul_In;
  input clock, reset, EnableChange;
  output we1, we2, we3, we4, WE, EOC_Flag, sig_OP;
  wire   FlagX, FlagY, DiagonalDoneX, DiagonalDoneY, WireX, WireY,
         DiagonalXDone, CompStart, EOF, \MainCount1[0] , signal, signal2, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903;
  wire   [10:0] Y_ramX;
  wire   [10:0] Y_ramY;
  wire   [255:0] RowX;
  wire   [255:0] RowY;
  wire   [10:0] Row_noX;
  wire   [10:0] Row_noY;
  wire   [1:0] FoundX;
  wire   [1:0] FoundY;
  wire   [255:0] NewRowX;
  wire   [255:0] NewRowY;
  wire   [12:0] PosDX;
  wire   [255:0] PaddedRow;
  wire   [47:0] NewDiagonalX;
  wire   [47:0] NewDiagonalY;
  wire   [47:0] ArbiterElement;
  wire   [12:0] ArbiterPos;
  wire   [255:0] OutputPaddedRow;
  wire   [12:0] PosDY;
  wire   [12:0] PosRowX;
  wire   [12:0] PosRowY;
  wire   [10:0] ComputeReq;
  wire   [255:0] OutputCompute;
  wire   [47:0] DiagonalX;
  wire   [47:0] DiagonalY;
  wire   [47:0] ElementUpdate;
  wire   [2:0] count;
  wire   [47:0] outA;
  wire   [48:0] outB;
  wire   [10:0] ElementAddr;
  wire   [47:0] d1;
  wire   [47:0] d2;
  wire   [47:0] d3;
  wire   [47:0] d4;
  wire   [47:0] d5;
  wire   [47:0] d6;
  wire   [47:0] d7;
  wire   [47:0] d8;
  wire   [47:0] d9;
  wire   [47:0] d10;
  wire   [47:0] d11;
  wire   [47:0] d12;
  wire   [47:0] d13;
  wire   [47:0] d14;
  wire   [47:0] d16;
  wire   [47:0] d17;
  wire   [24:0] adder_output;
  wire   [47:0] d18;
  wire   [48:0] SyncY;
  wire   [24:0] adder_output_imag;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4;

  DFF_X1 \d16_reg[47]  ( .D(subOut[47]), .CK(clock), .Q(d16[47]) );
  DFF_X1 \d17_reg[47]  ( .D(d16[47]), .CK(clock), .Q(d17[47]) );
  DFF_X1 \d18_reg[47]  ( .D(d17[47]), .CK(clock), .Q(d18[47]) );
  DFF_X1 \d16_reg[46]  ( .D(subOut[46]), .CK(clock), .Q(d16[46]) );
  DFF_X1 \d17_reg[46]  ( .D(d16[46]), .CK(clock), .Q(d17[46]) );
  DFF_X1 \d18_reg[46]  ( .D(d17[46]), .CK(clock), .Q(d18[46]) );
  DFF_X1 \d16_reg[45]  ( .D(subOut[45]), .CK(clock), .Q(d16[45]) );
  DFF_X1 \d17_reg[45]  ( .D(d16[45]), .CK(clock), .Q(d17[45]) );
  DFF_X1 \d18_reg[45]  ( .D(d17[45]), .CK(clock), .Q(d18[45]) );
  DFF_X1 \d16_reg[44]  ( .D(subOut[44]), .CK(clock), .Q(d16[44]) );
  DFF_X1 \d17_reg[44]  ( .D(d16[44]), .CK(clock), .Q(d17[44]) );
  DFF_X1 \d18_reg[44]  ( .D(d17[44]), .CK(clock), .Q(d18[44]) );
  DFF_X1 \d16_reg[43]  ( .D(subOut[43]), .CK(clock), .Q(d16[43]) );
  DFF_X1 \d17_reg[43]  ( .D(d16[43]), .CK(clock), .Q(d17[43]) );
  DFF_X1 \d18_reg[43]  ( .D(d17[43]), .CK(clock), .Q(d18[43]) );
  DFF_X1 \d16_reg[42]  ( .D(subOut[42]), .CK(clock), .Q(d16[42]) );
  DFF_X1 \d17_reg[42]  ( .D(d16[42]), .CK(clock), .Q(d17[42]) );
  DFF_X1 \d18_reg[42]  ( .D(d17[42]), .CK(clock), .Q(d18[42]) );
  DFF_X1 \d16_reg[41]  ( .D(subOut[41]), .CK(clock), .Q(d16[41]) );
  DFF_X1 \d17_reg[41]  ( .D(d16[41]), .CK(clock), .Q(d17[41]) );
  DFF_X1 \d18_reg[41]  ( .D(d17[41]), .CK(clock), .Q(d18[41]) );
  DFF_X1 \d16_reg[40]  ( .D(subOut[40]), .CK(clock), .Q(d16[40]) );
  DFF_X1 \d17_reg[40]  ( .D(d16[40]), .CK(clock), .Q(d17[40]) );
  DFF_X1 \d18_reg[40]  ( .D(d17[40]), .CK(clock), .Q(d18[40]) );
  DFF_X1 \d16_reg[39]  ( .D(subOut[39]), .CK(clock), .Q(d16[39]) );
  DFF_X1 \d17_reg[39]  ( .D(d16[39]), .CK(clock), .Q(d17[39]) );
  DFF_X1 \d18_reg[39]  ( .D(d17[39]), .CK(clock), .Q(d18[39]) );
  DFF_X1 \d16_reg[38]  ( .D(subOut[38]), .CK(clock), .Q(d16[38]) );
  DFF_X1 \d17_reg[38]  ( .D(d16[38]), .CK(clock), .Q(d17[38]) );
  DFF_X1 \d18_reg[38]  ( .D(d17[38]), .CK(clock), .Q(d18[38]) );
  DFF_X1 \d16_reg[37]  ( .D(subOut[37]), .CK(clock), .Q(d16[37]) );
  DFF_X1 \d17_reg[37]  ( .D(d16[37]), .CK(clock), .Q(d17[37]) );
  DFF_X1 \d18_reg[37]  ( .D(d17[37]), .CK(clock), .Q(d18[37]) );
  DFF_X1 \d16_reg[36]  ( .D(subOut[36]), .CK(clock), .Q(d16[36]) );
  DFF_X1 \d17_reg[36]  ( .D(d16[36]), .CK(clock), .Q(d17[36]) );
  DFF_X1 \d18_reg[36]  ( .D(d17[36]), .CK(clock), .Q(d18[36]) );
  DFF_X1 \d16_reg[35]  ( .D(subOut[35]), .CK(clock), .Q(d16[35]) );
  DFF_X1 \d17_reg[35]  ( .D(d16[35]), .CK(clock), .Q(d17[35]) );
  DFF_X1 \d18_reg[35]  ( .D(d17[35]), .CK(clock), .Q(d18[35]) );
  DFF_X1 \d16_reg[34]  ( .D(subOut[34]), .CK(clock), .Q(d16[34]) );
  DFF_X1 \d17_reg[34]  ( .D(d16[34]), .CK(clock), .Q(d17[34]) );
  DFF_X1 \d18_reg[34]  ( .D(d17[34]), .CK(clock), .Q(d18[34]) );
  DFF_X1 \d16_reg[33]  ( .D(subOut[33]), .CK(clock), .Q(d16[33]) );
  DFF_X1 \d17_reg[33]  ( .D(d16[33]), .CK(clock), .Q(d17[33]) );
  DFF_X1 \d18_reg[33]  ( .D(d17[33]), .CK(clock), .Q(d18[33]) );
  DFF_X1 \d16_reg[32]  ( .D(subOut[32]), .CK(clock), .Q(d16[32]) );
  DFF_X1 \d17_reg[32]  ( .D(d16[32]), .CK(clock), .Q(d17[32]) );
  DFF_X1 \d18_reg[32]  ( .D(d17[32]), .CK(clock), .Q(d18[32]) );
  DFF_X1 \d16_reg[31]  ( .D(subOut[31]), .CK(clock), .Q(d16[31]) );
  DFF_X1 \d17_reg[31]  ( .D(d16[31]), .CK(clock), .Q(d17[31]) );
  DFF_X1 \d18_reg[31]  ( .D(d17[31]), .CK(clock), .Q(d18[31]) );
  DFF_X1 \d16_reg[30]  ( .D(subOut[30]), .CK(clock), .Q(d16[30]) );
  DFF_X1 \d17_reg[30]  ( .D(d16[30]), .CK(clock), .Q(d17[30]) );
  DFF_X1 \d18_reg[30]  ( .D(d17[30]), .CK(clock), .Q(d18[30]) );
  DFF_X1 \d16_reg[29]  ( .D(subOut[29]), .CK(clock), .Q(d16[29]) );
  DFF_X1 \d17_reg[29]  ( .D(d16[29]), .CK(clock), .Q(d17[29]) );
  DFF_X1 \d18_reg[29]  ( .D(d17[29]), .CK(clock), .Q(d18[29]) );
  DFF_X1 \d16_reg[28]  ( .D(subOut[28]), .CK(clock), .Q(d16[28]) );
  DFF_X1 \d17_reg[28]  ( .D(d16[28]), .CK(clock), .Q(d17[28]) );
  DFF_X1 \d18_reg[28]  ( .D(d17[28]), .CK(clock), .Q(d18[28]) );
  DFF_X1 \d16_reg[27]  ( .D(subOut[27]), .CK(clock), .Q(d16[27]) );
  DFF_X1 \d17_reg[27]  ( .D(d16[27]), .CK(clock), .Q(d17[27]) );
  DFF_X1 \d18_reg[27]  ( .D(d17[27]), .CK(clock), .Q(d18[27]) );
  DFF_X1 \d16_reg[26]  ( .D(subOut[26]), .CK(clock), .Q(d16[26]) );
  DFF_X1 \d17_reg[26]  ( .D(d16[26]), .CK(clock), .Q(d17[26]) );
  DFF_X1 \d18_reg[26]  ( .D(d17[26]), .CK(clock), .Q(d18[26]) );
  DFF_X1 \d16_reg[25]  ( .D(subOut[25]), .CK(clock), .Q(d16[25]) );
  DFF_X1 \d17_reg[25]  ( .D(d16[25]), .CK(clock), .Q(d17[25]) );
  DFF_X1 \d18_reg[25]  ( .D(d17[25]), .CK(clock), .Q(d18[25]) );
  DFF_X1 \d16_reg[24]  ( .D(subOut[24]), .CK(clock), .Q(d16[24]) );
  DFF_X1 \d17_reg[24]  ( .D(d16[24]), .CK(clock), .Q(d17[24]) );
  DFF_X1 \d18_reg[24]  ( .D(d17[24]), .CK(clock), .Q(d18[24]) );
  DFF_X1 \d16_reg[23]  ( .D(subOut[23]), .CK(clock), .Q(d16[23]) );
  DFF_X1 \d17_reg[23]  ( .D(d16[23]), .CK(clock), .Q(d17[23]) );
  DFF_X1 \d18_reg[23]  ( .D(d17[23]), .CK(clock), .Q(d18[23]) );
  DFF_X1 \d16_reg[22]  ( .D(subOut[22]), .CK(clock), .Q(d16[22]) );
  DFF_X1 \d17_reg[22]  ( .D(d16[22]), .CK(clock), .Q(d17[22]) );
  DFF_X1 \d18_reg[22]  ( .D(d17[22]), .CK(clock), .Q(d18[22]) );
  DFF_X1 \d16_reg[21]  ( .D(subOut[21]), .CK(clock), .Q(d16[21]) );
  DFF_X1 \d17_reg[21]  ( .D(d16[21]), .CK(clock), .Q(d17[21]) );
  DFF_X1 \d18_reg[21]  ( .D(d17[21]), .CK(clock), .Q(d18[21]) );
  DFF_X1 \d16_reg[20]  ( .D(subOut[20]), .CK(clock), .Q(d16[20]) );
  DFF_X1 \d17_reg[20]  ( .D(d16[20]), .CK(clock), .Q(d17[20]) );
  DFF_X1 \d18_reg[20]  ( .D(d17[20]), .CK(clock), .Q(d18[20]) );
  DFF_X1 \d16_reg[19]  ( .D(subOut[19]), .CK(clock), .Q(d16[19]) );
  DFF_X1 \d17_reg[19]  ( .D(d16[19]), .CK(clock), .Q(d17[19]) );
  DFF_X1 \d18_reg[19]  ( .D(d17[19]), .CK(clock), .Q(d18[19]) );
  DFF_X1 \d16_reg[18]  ( .D(subOut[18]), .CK(clock), .Q(d16[18]) );
  DFF_X1 \d17_reg[18]  ( .D(d16[18]), .CK(clock), .Q(d17[18]) );
  DFF_X1 \d18_reg[18]  ( .D(d17[18]), .CK(clock), .Q(d18[18]) );
  DFF_X1 \d16_reg[17]  ( .D(subOut[17]), .CK(clock), .Q(d16[17]) );
  DFF_X1 \d17_reg[17]  ( .D(d16[17]), .CK(clock), .Q(d17[17]) );
  DFF_X1 \d18_reg[17]  ( .D(d17[17]), .CK(clock), .Q(d18[17]) );
  DFF_X1 \d16_reg[16]  ( .D(subOut[16]), .CK(clock), .Q(d16[16]) );
  DFF_X1 \d17_reg[16]  ( .D(d16[16]), .CK(clock), .Q(d17[16]) );
  DFF_X1 \d18_reg[16]  ( .D(d17[16]), .CK(clock), .Q(d18[16]) );
  DFF_X1 \d16_reg[15]  ( .D(subOut[15]), .CK(clock), .Q(d16[15]) );
  DFF_X1 \d17_reg[15]  ( .D(d16[15]), .CK(clock), .Q(d17[15]) );
  DFF_X1 \d18_reg[15]  ( .D(d17[15]), .CK(clock), .Q(d18[15]) );
  DFF_X1 \d16_reg[14]  ( .D(subOut[14]), .CK(clock), .Q(d16[14]) );
  DFF_X1 \d17_reg[14]  ( .D(d16[14]), .CK(clock), .Q(d17[14]) );
  DFF_X1 \d18_reg[14]  ( .D(d17[14]), .CK(clock), .Q(d18[14]) );
  DFF_X1 \d16_reg[13]  ( .D(subOut[13]), .CK(clock), .Q(d16[13]) );
  DFF_X1 \d17_reg[13]  ( .D(d16[13]), .CK(clock), .Q(d17[13]) );
  DFF_X1 \d18_reg[13]  ( .D(d17[13]), .CK(clock), .Q(d18[13]) );
  DFF_X1 \d16_reg[12]  ( .D(subOut[12]), .CK(clock), .Q(d16[12]) );
  DFF_X1 \d17_reg[12]  ( .D(d16[12]), .CK(clock), .Q(d17[12]) );
  DFF_X1 \d18_reg[12]  ( .D(d17[12]), .CK(clock), .Q(d18[12]) );
  DFF_X1 \d16_reg[11]  ( .D(subOut[11]), .CK(clock), .Q(d16[11]) );
  DFF_X1 \d17_reg[11]  ( .D(d16[11]), .CK(clock), .Q(d17[11]) );
  DFF_X1 \d18_reg[11]  ( .D(d17[11]), .CK(clock), .Q(d18[11]) );
  DFF_X1 \d16_reg[10]  ( .D(subOut[10]), .CK(clock), .Q(d16[10]) );
  DFF_X1 \d17_reg[10]  ( .D(d16[10]), .CK(clock), .Q(d17[10]) );
  DFF_X1 \d18_reg[10]  ( .D(d17[10]), .CK(clock), .Q(d18[10]) );
  DFF_X1 \d16_reg[9]  ( .D(subOut[9]), .CK(clock), .Q(d16[9]) );
  DFF_X1 \d17_reg[9]  ( .D(d16[9]), .CK(clock), .Q(d17[9]) );
  DFF_X1 \d18_reg[9]  ( .D(d17[9]), .CK(clock), .Q(d18[9]) );
  DFF_X1 \d16_reg[8]  ( .D(subOut[8]), .CK(clock), .Q(d16[8]) );
  DFF_X1 \d17_reg[8]  ( .D(d16[8]), .CK(clock), .Q(d17[8]) );
  DFF_X1 \d18_reg[8]  ( .D(d17[8]), .CK(clock), .Q(d18[8]) );
  DFF_X1 \d16_reg[7]  ( .D(subOut[7]), .CK(clock), .Q(d16[7]) );
  DFF_X1 \d17_reg[7]  ( .D(d16[7]), .CK(clock), .Q(d17[7]) );
  DFF_X1 \d18_reg[7]  ( .D(d17[7]), .CK(clock), .Q(d18[7]) );
  DFF_X1 \d16_reg[6]  ( .D(subOut[6]), .CK(clock), .Q(d16[6]) );
  DFF_X1 \d17_reg[6]  ( .D(d16[6]), .CK(clock), .Q(d17[6]) );
  DFF_X1 \d18_reg[6]  ( .D(d17[6]), .CK(clock), .Q(d18[6]) );
  DFF_X1 \d16_reg[5]  ( .D(subOut[5]), .CK(clock), .Q(d16[5]) );
  DFF_X1 \d17_reg[5]  ( .D(d16[5]), .CK(clock), .Q(d17[5]) );
  DFF_X1 \d18_reg[5]  ( .D(d17[5]), .CK(clock), .Q(d18[5]) );
  DFF_X1 \d16_reg[4]  ( .D(subOut[4]), .CK(clock), .Q(d16[4]) );
  DFF_X1 \d17_reg[4]  ( .D(d16[4]), .CK(clock), .Q(d17[4]) );
  DFF_X1 \d18_reg[4]  ( .D(d17[4]), .CK(clock), .Q(d18[4]) );
  DFF_X1 \d16_reg[3]  ( .D(subOut[3]), .CK(clock), .Q(d16[3]) );
  DFF_X1 \d17_reg[3]  ( .D(d16[3]), .CK(clock), .Q(d17[3]) );
  DFF_X1 \d18_reg[3]  ( .D(d17[3]), .CK(clock), .Q(d18[3]) );
  DFF_X1 \d16_reg[2]  ( .D(subOut[2]), .CK(clock), .Q(d16[2]) );
  DFF_X1 \d17_reg[2]  ( .D(d16[2]), .CK(clock), .Q(d17[2]) );
  DFF_X1 \d18_reg[2]  ( .D(d17[2]), .CK(clock), .Q(d18[2]) );
  DFF_X1 \d16_reg[1]  ( .D(subOut[1]), .CK(clock), .Q(d16[1]) );
  DFF_X1 \d17_reg[1]  ( .D(d16[1]), .CK(clock), .Q(d17[1]) );
  DFF_X1 \d18_reg[1]  ( .D(d17[1]), .CK(clock), .Q(d18[1]) );
  DFF_X1 \d16_reg[0]  ( .D(subOut[0]), .CK(clock), .Q(d16[0]) );
  DFF_X1 \d17_reg[0]  ( .D(d16[0]), .CK(clock), .Q(d17[0]) );
  DFF_X1 \d18_reg[0]  ( .D(d17[0]), .CK(clock), .Q(d18[0]) );
  DFF_X1 \d1_reg[47]  ( .D(outA[47]), .CK(clock), .Q(d1[47]) );
  DFF_X1 \d2_reg[47]  ( .D(d1[47]), .CK(clock), .Q(d2[47]) );
  DFF_X1 \d3_reg[47]  ( .D(d2[47]), .CK(clock), .Q(d3[47]) );
  DFF_X1 \d4_reg[47]  ( .D(d3[47]), .CK(clock), .Q(d4[47]) );
  DFF_X1 \d5_reg[47]  ( .D(d4[47]), .CK(clock), .Q(d5[47]) );
  DFF_X1 \d6_reg[47]  ( .D(d5[47]), .CK(clock), .Q(d6[47]) );
  DFF_X1 \d7_reg[47]  ( .D(d6[47]), .CK(clock), .Q(d7[47]) );
  DFF_X1 \d8_reg[47]  ( .D(d7[47]), .CK(clock), .Q(d8[47]) );
  DFF_X1 \d9_reg[47]  ( .D(d8[47]), .CK(clock), .Q(d9[47]) );
  DFF_X1 \d10_reg[47]  ( .D(d9[47]), .CK(clock), .Q(d10[47]) );
  DFF_X1 \d11_reg[47]  ( .D(d10[47]), .CK(clock), .Q(d11[47]) );
  DFF_X1 \d12_reg[47]  ( .D(d11[47]), .CK(clock), .Q(d12[47]) );
  DFF_X1 \d13_reg[47]  ( .D(d12[47]), .CK(clock), .Q(d13[47]) );
  DFF_X1 \d14_reg[47]  ( .D(d13[47]), .CK(clock), .Q(d14[47]) );
  DFF_X1 \d15_reg[47]  ( .D(d14[47]), .CK(clock), .QN(n96) );
  DFF_X1 \d1_reg[46]  ( .D(outA[46]), .CK(clock), .Q(d1[46]) );
  DFF_X1 \d2_reg[46]  ( .D(d1[46]), .CK(clock), .Q(d2[46]) );
  DFF_X1 \d3_reg[46]  ( .D(d2[46]), .CK(clock), .Q(d3[46]) );
  DFF_X1 \d4_reg[46]  ( .D(d3[46]), .CK(clock), .Q(d4[46]) );
  DFF_X1 \d5_reg[46]  ( .D(d4[46]), .CK(clock), .Q(d5[46]) );
  DFF_X1 \d6_reg[46]  ( .D(d5[46]), .CK(clock), .Q(d6[46]) );
  DFF_X1 \d7_reg[46]  ( .D(d6[46]), .CK(clock), .Q(d7[46]) );
  DFF_X1 \d8_reg[46]  ( .D(d7[46]), .CK(clock), .Q(d8[46]) );
  DFF_X1 \d9_reg[46]  ( .D(d8[46]), .CK(clock), .Q(d9[46]) );
  DFF_X1 \d10_reg[46]  ( .D(d9[46]), .CK(clock), .Q(d10[46]) );
  DFF_X1 \d11_reg[46]  ( .D(d10[46]), .CK(clock), .Q(d11[46]) );
  DFF_X1 \d12_reg[46]  ( .D(d11[46]), .CK(clock), .Q(d12[46]) );
  DFF_X1 \d13_reg[46]  ( .D(d12[46]), .CK(clock), .Q(d13[46]) );
  DFF_X1 \d14_reg[46]  ( .D(d13[46]), .CK(clock), .Q(d14[46]) );
  DFF_X1 \d15_reg[46]  ( .D(d14[46]), .CK(clock), .QN(n94) );
  DFF_X1 \d1_reg[45]  ( .D(outA[45]), .CK(clock), .Q(d1[45]) );
  DFF_X1 \d2_reg[45]  ( .D(d1[45]), .CK(clock), .Q(d2[45]) );
  DFF_X1 \d3_reg[45]  ( .D(d2[45]), .CK(clock), .Q(d3[45]) );
  DFF_X1 \d4_reg[45]  ( .D(d3[45]), .CK(clock), .Q(d4[45]) );
  DFF_X1 \d5_reg[45]  ( .D(d4[45]), .CK(clock), .Q(d5[45]) );
  DFF_X1 \d6_reg[45]  ( .D(d5[45]), .CK(clock), .Q(d6[45]) );
  DFF_X1 \d7_reg[45]  ( .D(d6[45]), .CK(clock), .Q(d7[45]) );
  DFF_X1 \d8_reg[45]  ( .D(d7[45]), .CK(clock), .Q(d8[45]) );
  DFF_X1 \d9_reg[45]  ( .D(d8[45]), .CK(clock), .Q(d9[45]) );
  DFF_X1 \d10_reg[45]  ( .D(d9[45]), .CK(clock), .Q(d10[45]) );
  DFF_X1 \d11_reg[45]  ( .D(d10[45]), .CK(clock), .Q(d11[45]) );
  DFF_X1 \d12_reg[45]  ( .D(d11[45]), .CK(clock), .Q(d12[45]) );
  DFF_X1 \d13_reg[45]  ( .D(d12[45]), .CK(clock), .Q(d13[45]) );
  DFF_X1 \d14_reg[45]  ( .D(d13[45]), .CK(clock), .Q(d14[45]) );
  DFF_X1 \d15_reg[45]  ( .D(d14[45]), .CK(clock), .QN(n92) );
  DFF_X1 \d1_reg[44]  ( .D(outA[44]), .CK(clock), .Q(d1[44]) );
  DFF_X1 \d2_reg[44]  ( .D(d1[44]), .CK(clock), .Q(d2[44]) );
  DFF_X1 \d3_reg[44]  ( .D(d2[44]), .CK(clock), .Q(d3[44]) );
  DFF_X1 \d4_reg[44]  ( .D(d3[44]), .CK(clock), .Q(d4[44]) );
  DFF_X1 \d5_reg[44]  ( .D(d4[44]), .CK(clock), .Q(d5[44]) );
  DFF_X1 \d6_reg[44]  ( .D(d5[44]), .CK(clock), .Q(d6[44]) );
  DFF_X1 \d7_reg[44]  ( .D(d6[44]), .CK(clock), .Q(d7[44]) );
  DFF_X1 \d8_reg[44]  ( .D(d7[44]), .CK(clock), .Q(d8[44]) );
  DFF_X1 \d9_reg[44]  ( .D(d8[44]), .CK(clock), .Q(d9[44]) );
  DFF_X1 \d10_reg[44]  ( .D(d9[44]), .CK(clock), .Q(d10[44]) );
  DFF_X1 \d11_reg[44]  ( .D(d10[44]), .CK(clock), .Q(d11[44]) );
  DFF_X1 \d12_reg[44]  ( .D(d11[44]), .CK(clock), .Q(d12[44]) );
  DFF_X1 \d13_reg[44]  ( .D(d12[44]), .CK(clock), .Q(d13[44]) );
  DFF_X1 \d14_reg[44]  ( .D(d13[44]), .CK(clock), .Q(d14[44]) );
  DFF_X1 \d15_reg[44]  ( .D(d14[44]), .CK(clock), .QN(n90) );
  DFF_X1 \d1_reg[43]  ( .D(outA[43]), .CK(clock), .Q(d1[43]) );
  DFF_X1 \d2_reg[43]  ( .D(d1[43]), .CK(clock), .Q(d2[43]) );
  DFF_X1 \d3_reg[43]  ( .D(d2[43]), .CK(clock), .Q(d3[43]) );
  DFF_X1 \d4_reg[43]  ( .D(d3[43]), .CK(clock), .Q(d4[43]) );
  DFF_X1 \d5_reg[43]  ( .D(d4[43]), .CK(clock), .Q(d5[43]) );
  DFF_X1 \d6_reg[43]  ( .D(d5[43]), .CK(clock), .Q(d6[43]) );
  DFF_X1 \d7_reg[43]  ( .D(d6[43]), .CK(clock), .Q(d7[43]) );
  DFF_X1 \d8_reg[43]  ( .D(d7[43]), .CK(clock), .Q(d8[43]) );
  DFF_X1 \d9_reg[43]  ( .D(d8[43]), .CK(clock), .Q(d9[43]) );
  DFF_X1 \d10_reg[43]  ( .D(d9[43]), .CK(clock), .Q(d10[43]) );
  DFF_X1 \d11_reg[43]  ( .D(d10[43]), .CK(clock), .Q(d11[43]) );
  DFF_X1 \d12_reg[43]  ( .D(d11[43]), .CK(clock), .Q(d12[43]) );
  DFF_X1 \d13_reg[43]  ( .D(d12[43]), .CK(clock), .Q(d13[43]) );
  DFF_X1 \d14_reg[43]  ( .D(d13[43]), .CK(clock), .Q(d14[43]) );
  DFF_X1 \d15_reg[43]  ( .D(d14[43]), .CK(clock), .QN(n88) );
  DFF_X1 \d1_reg[42]  ( .D(outA[42]), .CK(clock), .Q(d1[42]) );
  DFF_X1 \d2_reg[42]  ( .D(d1[42]), .CK(clock), .Q(d2[42]) );
  DFF_X1 \d3_reg[42]  ( .D(d2[42]), .CK(clock), .Q(d3[42]) );
  DFF_X1 \d4_reg[42]  ( .D(d3[42]), .CK(clock), .Q(d4[42]) );
  DFF_X1 \d5_reg[42]  ( .D(d4[42]), .CK(clock), .Q(d5[42]) );
  DFF_X1 \d6_reg[42]  ( .D(d5[42]), .CK(clock), .Q(d6[42]) );
  DFF_X1 \d7_reg[42]  ( .D(d6[42]), .CK(clock), .Q(d7[42]) );
  DFF_X1 \d8_reg[42]  ( .D(d7[42]), .CK(clock), .Q(d8[42]) );
  DFF_X1 \d9_reg[42]  ( .D(d8[42]), .CK(clock), .Q(d9[42]) );
  DFF_X1 \d10_reg[42]  ( .D(d9[42]), .CK(clock), .Q(d10[42]) );
  DFF_X1 \d11_reg[42]  ( .D(d10[42]), .CK(clock), .Q(d11[42]) );
  DFF_X1 \d12_reg[42]  ( .D(d11[42]), .CK(clock), .Q(d12[42]) );
  DFF_X1 \d13_reg[42]  ( .D(d12[42]), .CK(clock), .Q(d13[42]) );
  DFF_X1 \d14_reg[42]  ( .D(d13[42]), .CK(clock), .Q(d14[42]) );
  DFF_X1 \d15_reg[42]  ( .D(d14[42]), .CK(clock), .QN(n86) );
  DFF_X1 \d1_reg[41]  ( .D(outA[41]), .CK(clock), .Q(d1[41]) );
  DFF_X1 \d2_reg[41]  ( .D(d1[41]), .CK(clock), .Q(d2[41]) );
  DFF_X1 \d3_reg[41]  ( .D(d2[41]), .CK(clock), .Q(d3[41]) );
  DFF_X1 \d4_reg[41]  ( .D(d3[41]), .CK(clock), .Q(d4[41]) );
  DFF_X1 \d5_reg[41]  ( .D(d4[41]), .CK(clock), .Q(d5[41]) );
  DFF_X1 \d6_reg[41]  ( .D(d5[41]), .CK(clock), .Q(d6[41]) );
  DFF_X1 \d7_reg[41]  ( .D(d6[41]), .CK(clock), .Q(d7[41]) );
  DFF_X1 \d8_reg[41]  ( .D(d7[41]), .CK(clock), .Q(d8[41]) );
  DFF_X1 \d9_reg[41]  ( .D(d8[41]), .CK(clock), .Q(d9[41]) );
  DFF_X1 \d10_reg[41]  ( .D(d9[41]), .CK(clock), .Q(d10[41]) );
  DFF_X1 \d11_reg[41]  ( .D(d10[41]), .CK(clock), .Q(d11[41]) );
  DFF_X1 \d12_reg[41]  ( .D(d11[41]), .CK(clock), .Q(d12[41]) );
  DFF_X1 \d13_reg[41]  ( .D(d12[41]), .CK(clock), .Q(d13[41]) );
  DFF_X1 \d14_reg[41]  ( .D(d13[41]), .CK(clock), .Q(d14[41]) );
  DFF_X1 \d15_reg[41]  ( .D(d14[41]), .CK(clock), .QN(n84) );
  DFF_X1 \d1_reg[40]  ( .D(outA[40]), .CK(clock), .Q(d1[40]) );
  DFF_X1 \d2_reg[40]  ( .D(d1[40]), .CK(clock), .Q(d2[40]) );
  DFF_X1 \d3_reg[40]  ( .D(d2[40]), .CK(clock), .Q(d3[40]) );
  DFF_X1 \d4_reg[40]  ( .D(d3[40]), .CK(clock), .Q(d4[40]) );
  DFF_X1 \d5_reg[40]  ( .D(d4[40]), .CK(clock), .Q(d5[40]) );
  DFF_X1 \d6_reg[40]  ( .D(d5[40]), .CK(clock), .Q(d6[40]) );
  DFF_X1 \d7_reg[40]  ( .D(d6[40]), .CK(clock), .Q(d7[40]) );
  DFF_X1 \d8_reg[40]  ( .D(d7[40]), .CK(clock), .Q(d8[40]) );
  DFF_X1 \d9_reg[40]  ( .D(d8[40]), .CK(clock), .Q(d9[40]) );
  DFF_X1 \d10_reg[40]  ( .D(d9[40]), .CK(clock), .Q(d10[40]) );
  DFF_X1 \d11_reg[40]  ( .D(d10[40]), .CK(clock), .Q(d11[40]) );
  DFF_X1 \d12_reg[40]  ( .D(d11[40]), .CK(clock), .Q(d12[40]) );
  DFF_X1 \d13_reg[40]  ( .D(d12[40]), .CK(clock), .Q(d13[40]) );
  DFF_X1 \d14_reg[40]  ( .D(d13[40]), .CK(clock), .Q(d14[40]) );
  DFF_X1 \d15_reg[40]  ( .D(d14[40]), .CK(clock), .QN(n82) );
  DFF_X1 \d1_reg[39]  ( .D(outA[39]), .CK(clock), .Q(d1[39]) );
  DFF_X1 \d2_reg[39]  ( .D(d1[39]), .CK(clock), .Q(d2[39]) );
  DFF_X1 \d3_reg[39]  ( .D(d2[39]), .CK(clock), .Q(d3[39]) );
  DFF_X1 \d4_reg[39]  ( .D(d3[39]), .CK(clock), .Q(d4[39]) );
  DFF_X1 \d5_reg[39]  ( .D(d4[39]), .CK(clock), .Q(d5[39]) );
  DFF_X1 \d6_reg[39]  ( .D(d5[39]), .CK(clock), .Q(d6[39]) );
  DFF_X1 \d7_reg[39]  ( .D(d6[39]), .CK(clock), .Q(d7[39]) );
  DFF_X1 \d8_reg[39]  ( .D(d7[39]), .CK(clock), .Q(d8[39]) );
  DFF_X1 \d9_reg[39]  ( .D(d8[39]), .CK(clock), .Q(d9[39]) );
  DFF_X1 \d10_reg[39]  ( .D(d9[39]), .CK(clock), .Q(d10[39]) );
  DFF_X1 \d11_reg[39]  ( .D(d10[39]), .CK(clock), .Q(d11[39]) );
  DFF_X1 \d12_reg[39]  ( .D(d11[39]), .CK(clock), .Q(d12[39]) );
  DFF_X1 \d13_reg[39]  ( .D(d12[39]), .CK(clock), .Q(d13[39]) );
  DFF_X1 \d14_reg[39]  ( .D(d13[39]), .CK(clock), .Q(d14[39]) );
  DFF_X1 \d15_reg[39]  ( .D(d14[39]), .CK(clock), .QN(n80) );
  DFF_X1 \d1_reg[38]  ( .D(outA[38]), .CK(clock), .Q(d1[38]) );
  DFF_X1 \d2_reg[38]  ( .D(d1[38]), .CK(clock), .Q(d2[38]) );
  DFF_X1 \d3_reg[38]  ( .D(d2[38]), .CK(clock), .Q(d3[38]) );
  DFF_X1 \d4_reg[38]  ( .D(d3[38]), .CK(clock), .Q(d4[38]) );
  DFF_X1 \d5_reg[38]  ( .D(d4[38]), .CK(clock), .Q(d5[38]) );
  DFF_X1 \d6_reg[38]  ( .D(d5[38]), .CK(clock), .Q(d6[38]) );
  DFF_X1 \d7_reg[38]  ( .D(d6[38]), .CK(clock), .Q(d7[38]) );
  DFF_X1 \d8_reg[38]  ( .D(d7[38]), .CK(clock), .Q(d8[38]) );
  DFF_X1 \d9_reg[38]  ( .D(d8[38]), .CK(clock), .Q(d9[38]) );
  DFF_X1 \d10_reg[38]  ( .D(d9[38]), .CK(clock), .Q(d10[38]) );
  DFF_X1 \d11_reg[38]  ( .D(d10[38]), .CK(clock), .Q(d11[38]) );
  DFF_X1 \d12_reg[38]  ( .D(d11[38]), .CK(clock), .Q(d12[38]) );
  DFF_X1 \d13_reg[38]  ( .D(d12[38]), .CK(clock), .Q(d13[38]) );
  DFF_X1 \d14_reg[38]  ( .D(d13[38]), .CK(clock), .Q(d14[38]) );
  DFF_X1 \d15_reg[38]  ( .D(d14[38]), .CK(clock), .QN(n78) );
  DFF_X1 \d1_reg[37]  ( .D(outA[37]), .CK(clock), .Q(d1[37]) );
  DFF_X1 \d2_reg[37]  ( .D(d1[37]), .CK(clock), .Q(d2[37]) );
  DFF_X1 \d3_reg[37]  ( .D(d2[37]), .CK(clock), .Q(d3[37]) );
  DFF_X1 \d4_reg[37]  ( .D(d3[37]), .CK(clock), .Q(d4[37]) );
  DFF_X1 \d5_reg[37]  ( .D(d4[37]), .CK(clock), .Q(d5[37]) );
  DFF_X1 \d6_reg[37]  ( .D(d5[37]), .CK(clock), .Q(d6[37]) );
  DFF_X1 \d7_reg[37]  ( .D(d6[37]), .CK(clock), .Q(d7[37]) );
  DFF_X1 \d8_reg[37]  ( .D(d7[37]), .CK(clock), .Q(d8[37]) );
  DFF_X1 \d9_reg[37]  ( .D(d8[37]), .CK(clock), .Q(d9[37]) );
  DFF_X1 \d10_reg[37]  ( .D(d9[37]), .CK(clock), .Q(d10[37]) );
  DFF_X1 \d11_reg[37]  ( .D(d10[37]), .CK(clock), .Q(d11[37]) );
  DFF_X1 \d12_reg[37]  ( .D(d11[37]), .CK(clock), .Q(d12[37]) );
  DFF_X1 \d13_reg[37]  ( .D(d12[37]), .CK(clock), .Q(d13[37]) );
  DFF_X1 \d14_reg[37]  ( .D(d13[37]), .CK(clock), .Q(d14[37]) );
  DFF_X1 \d15_reg[37]  ( .D(d14[37]), .CK(clock), .QN(n76) );
  DFF_X1 \d1_reg[36]  ( .D(outA[36]), .CK(clock), .Q(d1[36]) );
  DFF_X1 \d2_reg[36]  ( .D(d1[36]), .CK(clock), .Q(d2[36]) );
  DFF_X1 \d3_reg[36]  ( .D(d2[36]), .CK(clock), .Q(d3[36]) );
  DFF_X1 \d4_reg[36]  ( .D(d3[36]), .CK(clock), .Q(d4[36]) );
  DFF_X1 \d5_reg[36]  ( .D(d4[36]), .CK(clock), .Q(d5[36]) );
  DFF_X1 \d6_reg[36]  ( .D(d5[36]), .CK(clock), .Q(d6[36]) );
  DFF_X1 \d7_reg[36]  ( .D(d6[36]), .CK(clock), .Q(d7[36]) );
  DFF_X1 \d8_reg[36]  ( .D(d7[36]), .CK(clock), .Q(d8[36]) );
  DFF_X1 \d9_reg[36]  ( .D(d8[36]), .CK(clock), .Q(d9[36]) );
  DFF_X1 \d10_reg[36]  ( .D(d9[36]), .CK(clock), .Q(d10[36]) );
  DFF_X1 \d11_reg[36]  ( .D(d10[36]), .CK(clock), .Q(d11[36]) );
  DFF_X1 \d12_reg[36]  ( .D(d11[36]), .CK(clock), .Q(d12[36]) );
  DFF_X1 \d13_reg[36]  ( .D(d12[36]), .CK(clock), .Q(d13[36]) );
  DFF_X1 \d14_reg[36]  ( .D(d13[36]), .CK(clock), .Q(d14[36]) );
  DFF_X1 \d15_reg[36]  ( .D(d14[36]), .CK(clock), .QN(n74) );
  DFF_X1 \d1_reg[35]  ( .D(outA[35]), .CK(clock), .Q(d1[35]) );
  DFF_X1 \d2_reg[35]  ( .D(d1[35]), .CK(clock), .Q(d2[35]) );
  DFF_X1 \d3_reg[35]  ( .D(d2[35]), .CK(clock), .Q(d3[35]) );
  DFF_X1 \d4_reg[35]  ( .D(d3[35]), .CK(clock), .Q(d4[35]) );
  DFF_X1 \d5_reg[35]  ( .D(d4[35]), .CK(clock), .Q(d5[35]) );
  DFF_X1 \d6_reg[35]  ( .D(d5[35]), .CK(clock), .Q(d6[35]) );
  DFF_X1 \d7_reg[35]  ( .D(d6[35]), .CK(clock), .Q(d7[35]) );
  DFF_X1 \d8_reg[35]  ( .D(d7[35]), .CK(clock), .Q(d8[35]) );
  DFF_X1 \d9_reg[35]  ( .D(d8[35]), .CK(clock), .Q(d9[35]) );
  DFF_X1 \d10_reg[35]  ( .D(d9[35]), .CK(clock), .Q(d10[35]) );
  DFF_X1 \d11_reg[35]  ( .D(d10[35]), .CK(clock), .Q(d11[35]) );
  DFF_X1 \d12_reg[35]  ( .D(d11[35]), .CK(clock), .Q(d12[35]) );
  DFF_X1 \d13_reg[35]  ( .D(d12[35]), .CK(clock), .Q(d13[35]) );
  DFF_X1 \d14_reg[35]  ( .D(d13[35]), .CK(clock), .Q(d14[35]) );
  DFF_X1 \d15_reg[35]  ( .D(d14[35]), .CK(clock), .QN(n72) );
  DFF_X1 \d1_reg[34]  ( .D(outA[34]), .CK(clock), .Q(d1[34]) );
  DFF_X1 \d2_reg[34]  ( .D(d1[34]), .CK(clock), .Q(d2[34]) );
  DFF_X1 \d3_reg[34]  ( .D(d2[34]), .CK(clock), .Q(d3[34]) );
  DFF_X1 \d4_reg[34]  ( .D(d3[34]), .CK(clock), .Q(d4[34]) );
  DFF_X1 \d5_reg[34]  ( .D(d4[34]), .CK(clock), .Q(d5[34]) );
  DFF_X1 \d6_reg[34]  ( .D(d5[34]), .CK(clock), .Q(d6[34]) );
  DFF_X1 \d7_reg[34]  ( .D(d6[34]), .CK(clock), .Q(d7[34]) );
  DFF_X1 \d8_reg[34]  ( .D(d7[34]), .CK(clock), .Q(d8[34]) );
  DFF_X1 \d9_reg[34]  ( .D(d8[34]), .CK(clock), .Q(d9[34]) );
  DFF_X1 \d10_reg[34]  ( .D(d9[34]), .CK(clock), .Q(d10[34]) );
  DFF_X1 \d11_reg[34]  ( .D(d10[34]), .CK(clock), .Q(d11[34]) );
  DFF_X1 \d12_reg[34]  ( .D(d11[34]), .CK(clock), .Q(d12[34]) );
  DFF_X1 \d13_reg[34]  ( .D(d12[34]), .CK(clock), .Q(d13[34]) );
  DFF_X1 \d14_reg[34]  ( .D(d13[34]), .CK(clock), .Q(d14[34]) );
  DFF_X1 \d15_reg[34]  ( .D(d14[34]), .CK(clock), .QN(n70) );
  DFF_X1 \d1_reg[33]  ( .D(outA[33]), .CK(clock), .Q(d1[33]) );
  DFF_X1 \d2_reg[33]  ( .D(d1[33]), .CK(clock), .Q(d2[33]) );
  DFF_X1 \d3_reg[33]  ( .D(d2[33]), .CK(clock), .Q(d3[33]) );
  DFF_X1 \d4_reg[33]  ( .D(d3[33]), .CK(clock), .Q(d4[33]) );
  DFF_X1 \d5_reg[33]  ( .D(d4[33]), .CK(clock), .Q(d5[33]) );
  DFF_X1 \d6_reg[33]  ( .D(d5[33]), .CK(clock), .Q(d6[33]) );
  DFF_X1 \d7_reg[33]  ( .D(d6[33]), .CK(clock), .Q(d7[33]) );
  DFF_X1 \d8_reg[33]  ( .D(d7[33]), .CK(clock), .Q(d8[33]) );
  DFF_X1 \d9_reg[33]  ( .D(d8[33]), .CK(clock), .Q(d9[33]) );
  DFF_X1 \d10_reg[33]  ( .D(d9[33]), .CK(clock), .Q(d10[33]) );
  DFF_X1 \d11_reg[33]  ( .D(d10[33]), .CK(clock), .Q(d11[33]) );
  DFF_X1 \d12_reg[33]  ( .D(d11[33]), .CK(clock), .Q(d12[33]) );
  DFF_X1 \d13_reg[33]  ( .D(d12[33]), .CK(clock), .Q(d13[33]) );
  DFF_X1 \d14_reg[33]  ( .D(d13[33]), .CK(clock), .Q(d14[33]) );
  DFF_X1 \d15_reg[33]  ( .D(d14[33]), .CK(clock), .QN(n68) );
  DFF_X1 \d1_reg[32]  ( .D(outA[32]), .CK(clock), .Q(d1[32]) );
  DFF_X1 \d2_reg[32]  ( .D(d1[32]), .CK(clock), .Q(d2[32]) );
  DFF_X1 \d3_reg[32]  ( .D(d2[32]), .CK(clock), .Q(d3[32]) );
  DFF_X1 \d4_reg[32]  ( .D(d3[32]), .CK(clock), .Q(d4[32]) );
  DFF_X1 \d5_reg[32]  ( .D(d4[32]), .CK(clock), .Q(d5[32]) );
  DFF_X1 \d6_reg[32]  ( .D(d5[32]), .CK(clock), .Q(d6[32]) );
  DFF_X1 \d7_reg[32]  ( .D(d6[32]), .CK(clock), .Q(d7[32]) );
  DFF_X1 \d8_reg[32]  ( .D(d7[32]), .CK(clock), .Q(d8[32]) );
  DFF_X1 \d9_reg[32]  ( .D(d8[32]), .CK(clock), .Q(d9[32]) );
  DFF_X1 \d10_reg[32]  ( .D(d9[32]), .CK(clock), .Q(d10[32]) );
  DFF_X1 \d11_reg[32]  ( .D(d10[32]), .CK(clock), .Q(d11[32]) );
  DFF_X1 \d12_reg[32]  ( .D(d11[32]), .CK(clock), .Q(d12[32]) );
  DFF_X1 \d13_reg[32]  ( .D(d12[32]), .CK(clock), .Q(d13[32]) );
  DFF_X1 \d14_reg[32]  ( .D(d13[32]), .CK(clock), .Q(d14[32]) );
  DFF_X1 \d15_reg[32]  ( .D(d14[32]), .CK(clock), .QN(n66) );
  DFF_X1 \d1_reg[31]  ( .D(outA[31]), .CK(clock), .Q(d1[31]) );
  DFF_X1 \d2_reg[31]  ( .D(d1[31]), .CK(clock), .Q(d2[31]) );
  DFF_X1 \d3_reg[31]  ( .D(d2[31]), .CK(clock), .Q(d3[31]) );
  DFF_X1 \d4_reg[31]  ( .D(d3[31]), .CK(clock), .Q(d4[31]) );
  DFF_X1 \d5_reg[31]  ( .D(d4[31]), .CK(clock), .Q(d5[31]) );
  DFF_X1 \d6_reg[31]  ( .D(d5[31]), .CK(clock), .Q(d6[31]) );
  DFF_X1 \d7_reg[31]  ( .D(d6[31]), .CK(clock), .Q(d7[31]) );
  DFF_X1 \d8_reg[31]  ( .D(d7[31]), .CK(clock), .Q(d8[31]) );
  DFF_X1 \d9_reg[31]  ( .D(d8[31]), .CK(clock), .Q(d9[31]) );
  DFF_X1 \d10_reg[31]  ( .D(d9[31]), .CK(clock), .Q(d10[31]) );
  DFF_X1 \d11_reg[31]  ( .D(d10[31]), .CK(clock), .Q(d11[31]) );
  DFF_X1 \d12_reg[31]  ( .D(d11[31]), .CK(clock), .Q(d12[31]) );
  DFF_X1 \d13_reg[31]  ( .D(d12[31]), .CK(clock), .Q(d13[31]) );
  DFF_X1 \d14_reg[31]  ( .D(d13[31]), .CK(clock), .Q(d14[31]) );
  DFF_X1 \d15_reg[31]  ( .D(d14[31]), .CK(clock), .QN(n64) );
  DFF_X1 \d1_reg[30]  ( .D(outA[30]), .CK(clock), .Q(d1[30]) );
  DFF_X1 \d2_reg[30]  ( .D(d1[30]), .CK(clock), .Q(d2[30]) );
  DFF_X1 \d3_reg[30]  ( .D(d2[30]), .CK(clock), .Q(d3[30]) );
  DFF_X1 \d4_reg[30]  ( .D(d3[30]), .CK(clock), .Q(d4[30]) );
  DFF_X1 \d5_reg[30]  ( .D(d4[30]), .CK(clock), .Q(d5[30]) );
  DFF_X1 \d6_reg[30]  ( .D(d5[30]), .CK(clock), .Q(d6[30]) );
  DFF_X1 \d7_reg[30]  ( .D(d6[30]), .CK(clock), .Q(d7[30]) );
  DFF_X1 \d8_reg[30]  ( .D(d7[30]), .CK(clock), .Q(d8[30]) );
  DFF_X1 \d9_reg[30]  ( .D(d8[30]), .CK(clock), .Q(d9[30]) );
  DFF_X1 \d10_reg[30]  ( .D(d9[30]), .CK(clock), .Q(d10[30]) );
  DFF_X1 \d11_reg[30]  ( .D(d10[30]), .CK(clock), .Q(d11[30]) );
  DFF_X1 \d12_reg[30]  ( .D(d11[30]), .CK(clock), .Q(d12[30]) );
  DFF_X1 \d13_reg[30]  ( .D(d12[30]), .CK(clock), .Q(d13[30]) );
  DFF_X1 \d14_reg[30]  ( .D(d13[30]), .CK(clock), .Q(d14[30]) );
  DFF_X1 \d15_reg[30]  ( .D(d14[30]), .CK(clock), .QN(n62) );
  DFF_X1 \d1_reg[29]  ( .D(outA[29]), .CK(clock), .Q(d1[29]) );
  DFF_X1 \d2_reg[29]  ( .D(d1[29]), .CK(clock), .Q(d2[29]) );
  DFF_X1 \d3_reg[29]  ( .D(d2[29]), .CK(clock), .Q(d3[29]) );
  DFF_X1 \d4_reg[29]  ( .D(d3[29]), .CK(clock), .Q(d4[29]) );
  DFF_X1 \d5_reg[29]  ( .D(d4[29]), .CK(clock), .Q(d5[29]) );
  DFF_X1 \d6_reg[29]  ( .D(d5[29]), .CK(clock), .Q(d6[29]) );
  DFF_X1 \d7_reg[29]  ( .D(d6[29]), .CK(clock), .Q(d7[29]) );
  DFF_X1 \d8_reg[29]  ( .D(d7[29]), .CK(clock), .Q(d8[29]) );
  DFF_X1 \d9_reg[29]  ( .D(d8[29]), .CK(clock), .Q(d9[29]) );
  DFF_X1 \d10_reg[29]  ( .D(d9[29]), .CK(clock), .Q(d10[29]) );
  DFF_X1 \d11_reg[29]  ( .D(d10[29]), .CK(clock), .Q(d11[29]) );
  DFF_X1 \d12_reg[29]  ( .D(d11[29]), .CK(clock), .Q(d12[29]) );
  DFF_X1 \d13_reg[29]  ( .D(d12[29]), .CK(clock), .Q(d13[29]) );
  DFF_X1 \d14_reg[29]  ( .D(d13[29]), .CK(clock), .Q(d14[29]) );
  DFF_X1 \d15_reg[29]  ( .D(d14[29]), .CK(clock), .QN(n60) );
  DFF_X1 \d1_reg[28]  ( .D(outA[28]), .CK(clock), .Q(d1[28]) );
  DFF_X1 \d2_reg[28]  ( .D(d1[28]), .CK(clock), .Q(d2[28]) );
  DFF_X1 \d3_reg[28]  ( .D(d2[28]), .CK(clock), .Q(d3[28]) );
  DFF_X1 \d4_reg[28]  ( .D(d3[28]), .CK(clock), .Q(d4[28]) );
  DFF_X1 \d5_reg[28]  ( .D(d4[28]), .CK(clock), .Q(d5[28]) );
  DFF_X1 \d6_reg[28]  ( .D(d5[28]), .CK(clock), .Q(d6[28]) );
  DFF_X1 \d7_reg[28]  ( .D(d6[28]), .CK(clock), .Q(d7[28]) );
  DFF_X1 \d8_reg[28]  ( .D(d7[28]), .CK(clock), .Q(d8[28]) );
  DFF_X1 \d9_reg[28]  ( .D(d8[28]), .CK(clock), .Q(d9[28]) );
  DFF_X1 \d10_reg[28]  ( .D(d9[28]), .CK(clock), .Q(d10[28]) );
  DFF_X1 \d11_reg[28]  ( .D(d10[28]), .CK(clock), .Q(d11[28]) );
  DFF_X1 \d12_reg[28]  ( .D(d11[28]), .CK(clock), .Q(d12[28]) );
  DFF_X1 \d13_reg[28]  ( .D(d12[28]), .CK(clock), .Q(d13[28]) );
  DFF_X1 \d14_reg[28]  ( .D(d13[28]), .CK(clock), .Q(d14[28]) );
  DFF_X1 \d15_reg[28]  ( .D(d14[28]), .CK(clock), .QN(n58) );
  DFF_X1 \d1_reg[27]  ( .D(outA[27]), .CK(clock), .Q(d1[27]) );
  DFF_X1 \d2_reg[27]  ( .D(d1[27]), .CK(clock), .Q(d2[27]) );
  DFF_X1 \d3_reg[27]  ( .D(d2[27]), .CK(clock), .Q(d3[27]) );
  DFF_X1 \d4_reg[27]  ( .D(d3[27]), .CK(clock), .Q(d4[27]) );
  DFF_X1 \d5_reg[27]  ( .D(d4[27]), .CK(clock), .Q(d5[27]) );
  DFF_X1 \d6_reg[27]  ( .D(d5[27]), .CK(clock), .Q(d6[27]) );
  DFF_X1 \d7_reg[27]  ( .D(d6[27]), .CK(clock), .Q(d7[27]) );
  DFF_X1 \d8_reg[27]  ( .D(d7[27]), .CK(clock), .Q(d8[27]) );
  DFF_X1 \d9_reg[27]  ( .D(d8[27]), .CK(clock), .Q(d9[27]) );
  DFF_X1 \d10_reg[27]  ( .D(d9[27]), .CK(clock), .Q(d10[27]) );
  DFF_X1 \d11_reg[27]  ( .D(d10[27]), .CK(clock), .Q(d11[27]) );
  DFF_X1 \d12_reg[27]  ( .D(d11[27]), .CK(clock), .Q(d12[27]) );
  DFF_X1 \d13_reg[27]  ( .D(d12[27]), .CK(clock), .Q(d13[27]) );
  DFF_X1 \d14_reg[27]  ( .D(d13[27]), .CK(clock), .Q(d14[27]) );
  DFF_X1 \d15_reg[27]  ( .D(d14[27]), .CK(clock), .QN(n56) );
  DFF_X1 \d1_reg[26]  ( .D(outA[26]), .CK(clock), .Q(d1[26]) );
  DFF_X1 \d2_reg[26]  ( .D(d1[26]), .CK(clock), .Q(d2[26]) );
  DFF_X1 \d3_reg[26]  ( .D(d2[26]), .CK(clock), .Q(d3[26]) );
  DFF_X1 \d4_reg[26]  ( .D(d3[26]), .CK(clock), .Q(d4[26]) );
  DFF_X1 \d5_reg[26]  ( .D(d4[26]), .CK(clock), .Q(d5[26]) );
  DFF_X1 \d6_reg[26]  ( .D(d5[26]), .CK(clock), .Q(d6[26]) );
  DFF_X1 \d7_reg[26]  ( .D(d6[26]), .CK(clock), .Q(d7[26]) );
  DFF_X1 \d8_reg[26]  ( .D(d7[26]), .CK(clock), .Q(d8[26]) );
  DFF_X1 \d9_reg[26]  ( .D(d8[26]), .CK(clock), .Q(d9[26]) );
  DFF_X1 \d10_reg[26]  ( .D(d9[26]), .CK(clock), .Q(d10[26]) );
  DFF_X1 \d11_reg[26]  ( .D(d10[26]), .CK(clock), .Q(d11[26]) );
  DFF_X1 \d12_reg[26]  ( .D(d11[26]), .CK(clock), .Q(d12[26]) );
  DFF_X1 \d13_reg[26]  ( .D(d12[26]), .CK(clock), .Q(d13[26]) );
  DFF_X1 \d14_reg[26]  ( .D(d13[26]), .CK(clock), .Q(d14[26]) );
  DFF_X1 \d15_reg[26]  ( .D(d14[26]), .CK(clock), .QN(n54) );
  DFF_X1 \d1_reg[25]  ( .D(outA[25]), .CK(clock), .Q(d1[25]) );
  DFF_X1 \d2_reg[25]  ( .D(d1[25]), .CK(clock), .Q(d2[25]) );
  DFF_X1 \d3_reg[25]  ( .D(d2[25]), .CK(clock), .Q(d3[25]) );
  DFF_X1 \d4_reg[25]  ( .D(d3[25]), .CK(clock), .Q(d4[25]) );
  DFF_X1 \d5_reg[25]  ( .D(d4[25]), .CK(clock), .Q(d5[25]) );
  DFF_X1 \d6_reg[25]  ( .D(d5[25]), .CK(clock), .Q(d6[25]) );
  DFF_X1 \d7_reg[25]  ( .D(d6[25]), .CK(clock), .Q(d7[25]) );
  DFF_X1 \d8_reg[25]  ( .D(d7[25]), .CK(clock), .Q(d8[25]) );
  DFF_X1 \d9_reg[25]  ( .D(d8[25]), .CK(clock), .Q(d9[25]) );
  DFF_X1 \d10_reg[25]  ( .D(d9[25]), .CK(clock), .Q(d10[25]) );
  DFF_X1 \d11_reg[25]  ( .D(d10[25]), .CK(clock), .Q(d11[25]) );
  DFF_X1 \d12_reg[25]  ( .D(d11[25]), .CK(clock), .Q(d12[25]) );
  DFF_X1 \d13_reg[25]  ( .D(d12[25]), .CK(clock), .Q(d13[25]) );
  DFF_X1 \d14_reg[25]  ( .D(d13[25]), .CK(clock), .Q(d14[25]) );
  DFF_X1 \d15_reg[25]  ( .D(d14[25]), .CK(clock), .QN(n52) );
  DFF_X1 \d1_reg[24]  ( .D(outA[24]), .CK(clock), .Q(d1[24]) );
  DFF_X1 \d2_reg[24]  ( .D(d1[24]), .CK(clock), .Q(d2[24]) );
  DFF_X1 \d3_reg[24]  ( .D(d2[24]), .CK(clock), .Q(d3[24]) );
  DFF_X1 \d4_reg[24]  ( .D(d3[24]), .CK(clock), .Q(d4[24]) );
  DFF_X1 \d5_reg[24]  ( .D(d4[24]), .CK(clock), .Q(d5[24]) );
  DFF_X1 \d6_reg[24]  ( .D(d5[24]), .CK(clock), .Q(d6[24]) );
  DFF_X1 \d7_reg[24]  ( .D(d6[24]), .CK(clock), .Q(d7[24]) );
  DFF_X1 \d8_reg[24]  ( .D(d7[24]), .CK(clock), .Q(d8[24]) );
  DFF_X1 \d9_reg[24]  ( .D(d8[24]), .CK(clock), .Q(d9[24]) );
  DFF_X1 \d10_reg[24]  ( .D(d9[24]), .CK(clock), .Q(d10[24]) );
  DFF_X1 \d11_reg[24]  ( .D(d10[24]), .CK(clock), .Q(d11[24]) );
  DFF_X1 \d12_reg[24]  ( .D(d11[24]), .CK(clock), .Q(d12[24]) );
  DFF_X1 \d13_reg[24]  ( .D(d12[24]), .CK(clock), .Q(d13[24]) );
  DFF_X1 \d14_reg[24]  ( .D(d13[24]), .CK(clock), .Q(d14[24]) );
  DFF_X1 \d15_reg[24]  ( .D(d14[24]), .CK(clock), .QN(n50) );
  DFF_X1 \d1_reg[23]  ( .D(outA[23]), .CK(clock), .Q(d1[23]) );
  DFF_X1 \d2_reg[23]  ( .D(d1[23]), .CK(clock), .Q(d2[23]) );
  DFF_X1 \d3_reg[23]  ( .D(d2[23]), .CK(clock), .Q(d3[23]) );
  DFF_X1 \d4_reg[23]  ( .D(d3[23]), .CK(clock), .Q(d4[23]) );
  DFF_X1 \d5_reg[23]  ( .D(d4[23]), .CK(clock), .Q(d5[23]) );
  DFF_X1 \d6_reg[23]  ( .D(d5[23]), .CK(clock), .Q(d6[23]) );
  DFF_X1 \d7_reg[23]  ( .D(d6[23]), .CK(clock), .Q(d7[23]) );
  DFF_X1 \d8_reg[23]  ( .D(d7[23]), .CK(clock), .Q(d8[23]) );
  DFF_X1 \d9_reg[23]  ( .D(d8[23]), .CK(clock), .Q(d9[23]) );
  DFF_X1 \d10_reg[23]  ( .D(d9[23]), .CK(clock), .Q(d10[23]) );
  DFF_X1 \d11_reg[23]  ( .D(d10[23]), .CK(clock), .Q(d11[23]) );
  DFF_X1 \d12_reg[23]  ( .D(d11[23]), .CK(clock), .Q(d12[23]) );
  DFF_X1 \d13_reg[23]  ( .D(d12[23]), .CK(clock), .Q(d13[23]) );
  DFF_X1 \d14_reg[23]  ( .D(d13[23]), .CK(clock), .Q(d14[23]) );
  DFF_X1 \d15_reg[23]  ( .D(d14[23]), .CK(clock), .QN(n48) );
  DFF_X1 \d1_reg[22]  ( .D(outA[22]), .CK(clock), .Q(d1[22]) );
  DFF_X1 \d2_reg[22]  ( .D(d1[22]), .CK(clock), .Q(d2[22]) );
  DFF_X1 \d3_reg[22]  ( .D(d2[22]), .CK(clock), .Q(d3[22]) );
  DFF_X1 \d4_reg[22]  ( .D(d3[22]), .CK(clock), .Q(d4[22]) );
  DFF_X1 \d5_reg[22]  ( .D(d4[22]), .CK(clock), .Q(d5[22]) );
  DFF_X1 \d6_reg[22]  ( .D(d5[22]), .CK(clock), .Q(d6[22]) );
  DFF_X1 \d7_reg[22]  ( .D(d6[22]), .CK(clock), .Q(d7[22]) );
  DFF_X1 \d8_reg[22]  ( .D(d7[22]), .CK(clock), .Q(d8[22]) );
  DFF_X1 \d9_reg[22]  ( .D(d8[22]), .CK(clock), .Q(d9[22]) );
  DFF_X1 \d10_reg[22]  ( .D(d9[22]), .CK(clock), .Q(d10[22]) );
  DFF_X1 \d11_reg[22]  ( .D(d10[22]), .CK(clock), .Q(d11[22]) );
  DFF_X1 \d12_reg[22]  ( .D(d11[22]), .CK(clock), .Q(d12[22]) );
  DFF_X1 \d13_reg[22]  ( .D(d12[22]), .CK(clock), .Q(d13[22]) );
  DFF_X1 \d14_reg[22]  ( .D(d13[22]), .CK(clock), .Q(d14[22]) );
  DFF_X1 \d15_reg[22]  ( .D(d14[22]), .CK(clock), .QN(n46) );
  DFF_X1 \d1_reg[21]  ( .D(outA[21]), .CK(clock), .Q(d1[21]) );
  DFF_X1 \d2_reg[21]  ( .D(d1[21]), .CK(clock), .Q(d2[21]) );
  DFF_X1 \d3_reg[21]  ( .D(d2[21]), .CK(clock), .Q(d3[21]) );
  DFF_X1 \d4_reg[21]  ( .D(d3[21]), .CK(clock), .Q(d4[21]) );
  DFF_X1 \d5_reg[21]  ( .D(d4[21]), .CK(clock), .Q(d5[21]) );
  DFF_X1 \d6_reg[21]  ( .D(d5[21]), .CK(clock), .Q(d6[21]) );
  DFF_X1 \d7_reg[21]  ( .D(d6[21]), .CK(clock), .Q(d7[21]) );
  DFF_X1 \d8_reg[21]  ( .D(d7[21]), .CK(clock), .Q(d8[21]) );
  DFF_X1 \d9_reg[21]  ( .D(d8[21]), .CK(clock), .Q(d9[21]) );
  DFF_X1 \d10_reg[21]  ( .D(d9[21]), .CK(clock), .Q(d10[21]) );
  DFF_X1 \d11_reg[21]  ( .D(d10[21]), .CK(clock), .Q(d11[21]) );
  DFF_X1 \d12_reg[21]  ( .D(d11[21]), .CK(clock), .Q(d12[21]) );
  DFF_X1 \d13_reg[21]  ( .D(d12[21]), .CK(clock), .Q(d13[21]) );
  DFF_X1 \d14_reg[21]  ( .D(d13[21]), .CK(clock), .Q(d14[21]) );
  DFF_X1 \d15_reg[21]  ( .D(d14[21]), .CK(clock), .QN(n44) );
  DFF_X1 \d1_reg[20]  ( .D(outA[20]), .CK(clock), .Q(d1[20]) );
  DFF_X1 \d2_reg[20]  ( .D(d1[20]), .CK(clock), .Q(d2[20]) );
  DFF_X1 \d3_reg[20]  ( .D(d2[20]), .CK(clock), .Q(d3[20]) );
  DFF_X1 \d4_reg[20]  ( .D(d3[20]), .CK(clock), .Q(d4[20]) );
  DFF_X1 \d5_reg[20]  ( .D(d4[20]), .CK(clock), .Q(d5[20]) );
  DFF_X1 \d6_reg[20]  ( .D(d5[20]), .CK(clock), .Q(d6[20]) );
  DFF_X1 \d7_reg[20]  ( .D(d6[20]), .CK(clock), .Q(d7[20]) );
  DFF_X1 \d8_reg[20]  ( .D(d7[20]), .CK(clock), .Q(d8[20]) );
  DFF_X1 \d9_reg[20]  ( .D(d8[20]), .CK(clock), .Q(d9[20]) );
  DFF_X1 \d10_reg[20]  ( .D(d9[20]), .CK(clock), .Q(d10[20]) );
  DFF_X1 \d11_reg[20]  ( .D(d10[20]), .CK(clock), .Q(d11[20]) );
  DFF_X1 \d12_reg[20]  ( .D(d11[20]), .CK(clock), .Q(d12[20]) );
  DFF_X1 \d13_reg[20]  ( .D(d12[20]), .CK(clock), .Q(d13[20]) );
  DFF_X1 \d14_reg[20]  ( .D(d13[20]), .CK(clock), .Q(d14[20]) );
  DFF_X1 \d15_reg[20]  ( .D(d14[20]), .CK(clock), .QN(n42) );
  DFF_X1 \d1_reg[19]  ( .D(outA[19]), .CK(clock), .Q(d1[19]) );
  DFF_X1 \d2_reg[19]  ( .D(d1[19]), .CK(clock), .Q(d2[19]) );
  DFF_X1 \d3_reg[19]  ( .D(d2[19]), .CK(clock), .Q(d3[19]) );
  DFF_X1 \d4_reg[19]  ( .D(d3[19]), .CK(clock), .Q(d4[19]) );
  DFF_X1 \d5_reg[19]  ( .D(d4[19]), .CK(clock), .Q(d5[19]) );
  DFF_X1 \d6_reg[19]  ( .D(d5[19]), .CK(clock), .Q(d6[19]) );
  DFF_X1 \d7_reg[19]  ( .D(d6[19]), .CK(clock), .Q(d7[19]) );
  DFF_X1 \d8_reg[19]  ( .D(d7[19]), .CK(clock), .Q(d8[19]) );
  DFF_X1 \d9_reg[19]  ( .D(d8[19]), .CK(clock), .Q(d9[19]) );
  DFF_X1 \d10_reg[19]  ( .D(d9[19]), .CK(clock), .Q(d10[19]) );
  DFF_X1 \d11_reg[19]  ( .D(d10[19]), .CK(clock), .Q(d11[19]) );
  DFF_X1 \d12_reg[19]  ( .D(d11[19]), .CK(clock), .Q(d12[19]) );
  DFF_X1 \d13_reg[19]  ( .D(d12[19]), .CK(clock), .Q(d13[19]) );
  DFF_X1 \d14_reg[19]  ( .D(d13[19]), .CK(clock), .Q(d14[19]) );
  DFF_X1 \d15_reg[19]  ( .D(d14[19]), .CK(clock), .QN(n40) );
  DFF_X1 \d1_reg[18]  ( .D(outA[18]), .CK(clock), .Q(d1[18]) );
  DFF_X1 \d2_reg[18]  ( .D(d1[18]), .CK(clock), .Q(d2[18]) );
  DFF_X1 \d3_reg[18]  ( .D(d2[18]), .CK(clock), .Q(d3[18]) );
  DFF_X1 \d4_reg[18]  ( .D(d3[18]), .CK(clock), .Q(d4[18]) );
  DFF_X1 \d5_reg[18]  ( .D(d4[18]), .CK(clock), .Q(d5[18]) );
  DFF_X1 \d6_reg[18]  ( .D(d5[18]), .CK(clock), .Q(d6[18]) );
  DFF_X1 \d7_reg[18]  ( .D(d6[18]), .CK(clock), .Q(d7[18]) );
  DFF_X1 \d8_reg[18]  ( .D(d7[18]), .CK(clock), .Q(d8[18]) );
  DFF_X1 \d9_reg[18]  ( .D(d8[18]), .CK(clock), .Q(d9[18]) );
  DFF_X1 \d10_reg[18]  ( .D(d9[18]), .CK(clock), .Q(d10[18]) );
  DFF_X1 \d11_reg[18]  ( .D(d10[18]), .CK(clock), .Q(d11[18]) );
  DFF_X1 \d12_reg[18]  ( .D(d11[18]), .CK(clock), .Q(d12[18]) );
  DFF_X1 \d13_reg[18]  ( .D(d12[18]), .CK(clock), .Q(d13[18]) );
  DFF_X1 \d14_reg[18]  ( .D(d13[18]), .CK(clock), .Q(d14[18]) );
  DFF_X1 \d15_reg[18]  ( .D(d14[18]), .CK(clock), .QN(n38) );
  DFF_X1 \d1_reg[17]  ( .D(outA[17]), .CK(clock), .Q(d1[17]) );
  DFF_X1 \d2_reg[17]  ( .D(d1[17]), .CK(clock), .Q(d2[17]) );
  DFF_X1 \d3_reg[17]  ( .D(d2[17]), .CK(clock), .Q(d3[17]) );
  DFF_X1 \d4_reg[17]  ( .D(d3[17]), .CK(clock), .Q(d4[17]) );
  DFF_X1 \d5_reg[17]  ( .D(d4[17]), .CK(clock), .Q(d5[17]) );
  DFF_X1 \d6_reg[17]  ( .D(d5[17]), .CK(clock), .Q(d6[17]) );
  DFF_X1 \d7_reg[17]  ( .D(d6[17]), .CK(clock), .Q(d7[17]) );
  DFF_X1 \d8_reg[17]  ( .D(d7[17]), .CK(clock), .Q(d8[17]) );
  DFF_X1 \d9_reg[17]  ( .D(d8[17]), .CK(clock), .Q(d9[17]) );
  DFF_X1 \d10_reg[17]  ( .D(d9[17]), .CK(clock), .Q(d10[17]) );
  DFF_X1 \d11_reg[17]  ( .D(d10[17]), .CK(clock), .Q(d11[17]) );
  DFF_X1 \d12_reg[17]  ( .D(d11[17]), .CK(clock), .Q(d12[17]) );
  DFF_X1 \d13_reg[17]  ( .D(d12[17]), .CK(clock), .Q(d13[17]) );
  DFF_X1 \d14_reg[17]  ( .D(d13[17]), .CK(clock), .Q(d14[17]) );
  DFF_X1 \d15_reg[17]  ( .D(d14[17]), .CK(clock), .QN(n36) );
  DFF_X1 \d1_reg[16]  ( .D(outA[16]), .CK(clock), .Q(d1[16]) );
  DFF_X1 \d2_reg[16]  ( .D(d1[16]), .CK(clock), .Q(d2[16]) );
  DFF_X1 \d3_reg[16]  ( .D(d2[16]), .CK(clock), .Q(d3[16]) );
  DFF_X1 \d4_reg[16]  ( .D(d3[16]), .CK(clock), .Q(d4[16]) );
  DFF_X1 \d5_reg[16]  ( .D(d4[16]), .CK(clock), .Q(d5[16]) );
  DFF_X1 \d6_reg[16]  ( .D(d5[16]), .CK(clock), .Q(d6[16]) );
  DFF_X1 \d7_reg[16]  ( .D(d6[16]), .CK(clock), .Q(d7[16]) );
  DFF_X1 \d8_reg[16]  ( .D(d7[16]), .CK(clock), .Q(d8[16]) );
  DFF_X1 \d9_reg[16]  ( .D(d8[16]), .CK(clock), .Q(d9[16]) );
  DFF_X1 \d10_reg[16]  ( .D(d9[16]), .CK(clock), .Q(d10[16]) );
  DFF_X1 \d11_reg[16]  ( .D(d10[16]), .CK(clock), .Q(d11[16]) );
  DFF_X1 \d12_reg[16]  ( .D(d11[16]), .CK(clock), .Q(d12[16]) );
  DFF_X1 \d13_reg[16]  ( .D(d12[16]), .CK(clock), .Q(d13[16]) );
  DFF_X1 \d14_reg[16]  ( .D(d13[16]), .CK(clock), .Q(d14[16]) );
  DFF_X1 \d15_reg[16]  ( .D(d14[16]), .CK(clock), .QN(n34) );
  DFF_X1 \d1_reg[15]  ( .D(outA[15]), .CK(clock), .Q(d1[15]) );
  DFF_X1 \d2_reg[15]  ( .D(d1[15]), .CK(clock), .Q(d2[15]) );
  DFF_X1 \d3_reg[15]  ( .D(d2[15]), .CK(clock), .Q(d3[15]) );
  DFF_X1 \d4_reg[15]  ( .D(d3[15]), .CK(clock), .Q(d4[15]) );
  DFF_X1 \d5_reg[15]  ( .D(d4[15]), .CK(clock), .Q(d5[15]) );
  DFF_X1 \d6_reg[15]  ( .D(d5[15]), .CK(clock), .Q(d6[15]) );
  DFF_X1 \d7_reg[15]  ( .D(d6[15]), .CK(clock), .Q(d7[15]) );
  DFF_X1 \d8_reg[15]  ( .D(d7[15]), .CK(clock), .Q(d8[15]) );
  DFF_X1 \d9_reg[15]  ( .D(d8[15]), .CK(clock), .Q(d9[15]) );
  DFF_X1 \d10_reg[15]  ( .D(d9[15]), .CK(clock), .Q(d10[15]) );
  DFF_X1 \d11_reg[15]  ( .D(d10[15]), .CK(clock), .Q(d11[15]) );
  DFF_X1 \d12_reg[15]  ( .D(d11[15]), .CK(clock), .Q(d12[15]) );
  DFF_X1 \d13_reg[15]  ( .D(d12[15]), .CK(clock), .Q(d13[15]) );
  DFF_X1 \d14_reg[15]  ( .D(d13[15]), .CK(clock), .Q(d14[15]) );
  DFF_X1 \d15_reg[15]  ( .D(d14[15]), .CK(clock), .QN(n32) );
  DFF_X1 \d1_reg[14]  ( .D(outA[14]), .CK(clock), .Q(d1[14]) );
  DFF_X1 \d2_reg[14]  ( .D(d1[14]), .CK(clock), .Q(d2[14]) );
  DFF_X1 \d3_reg[14]  ( .D(d2[14]), .CK(clock), .Q(d3[14]) );
  DFF_X1 \d4_reg[14]  ( .D(d3[14]), .CK(clock), .Q(d4[14]) );
  DFF_X1 \d5_reg[14]  ( .D(d4[14]), .CK(clock), .Q(d5[14]) );
  DFF_X1 \d6_reg[14]  ( .D(d5[14]), .CK(clock), .Q(d6[14]) );
  DFF_X1 \d7_reg[14]  ( .D(d6[14]), .CK(clock), .Q(d7[14]) );
  DFF_X1 \d8_reg[14]  ( .D(d7[14]), .CK(clock), .Q(d8[14]) );
  DFF_X1 \d9_reg[14]  ( .D(d8[14]), .CK(clock), .Q(d9[14]) );
  DFF_X1 \d10_reg[14]  ( .D(d9[14]), .CK(clock), .Q(d10[14]) );
  DFF_X1 \d11_reg[14]  ( .D(d10[14]), .CK(clock), .Q(d11[14]) );
  DFF_X1 \d12_reg[14]  ( .D(d11[14]), .CK(clock), .Q(d12[14]) );
  DFF_X1 \d13_reg[14]  ( .D(d12[14]), .CK(clock), .Q(d13[14]) );
  DFF_X1 \d14_reg[14]  ( .D(d13[14]), .CK(clock), .Q(d14[14]) );
  DFF_X1 \d15_reg[14]  ( .D(d14[14]), .CK(clock), .QN(n30) );
  DFF_X1 \d1_reg[13]  ( .D(outA[13]), .CK(clock), .Q(d1[13]) );
  DFF_X1 \d2_reg[13]  ( .D(d1[13]), .CK(clock), .Q(d2[13]) );
  DFF_X1 \d3_reg[13]  ( .D(d2[13]), .CK(clock), .Q(d3[13]) );
  DFF_X1 \d4_reg[13]  ( .D(d3[13]), .CK(clock), .Q(d4[13]) );
  DFF_X1 \d5_reg[13]  ( .D(d4[13]), .CK(clock), .Q(d5[13]) );
  DFF_X1 \d6_reg[13]  ( .D(d5[13]), .CK(clock), .Q(d6[13]) );
  DFF_X1 \d7_reg[13]  ( .D(d6[13]), .CK(clock), .Q(d7[13]) );
  DFF_X1 \d8_reg[13]  ( .D(d7[13]), .CK(clock), .Q(d8[13]) );
  DFF_X1 \d9_reg[13]  ( .D(d8[13]), .CK(clock), .Q(d9[13]) );
  DFF_X1 \d10_reg[13]  ( .D(d9[13]), .CK(clock), .Q(d10[13]) );
  DFF_X1 \d11_reg[13]  ( .D(d10[13]), .CK(clock), .Q(d11[13]) );
  DFF_X1 \d12_reg[13]  ( .D(d11[13]), .CK(clock), .Q(d12[13]) );
  DFF_X1 \d13_reg[13]  ( .D(d12[13]), .CK(clock), .Q(d13[13]) );
  DFF_X1 \d14_reg[13]  ( .D(d13[13]), .CK(clock), .Q(d14[13]) );
  DFF_X1 \d15_reg[13]  ( .D(d14[13]), .CK(clock), .QN(n28) );
  DFF_X1 \d1_reg[12]  ( .D(outA[12]), .CK(clock), .Q(d1[12]) );
  DFF_X1 \d2_reg[12]  ( .D(d1[12]), .CK(clock), .Q(d2[12]) );
  DFF_X1 \d3_reg[12]  ( .D(d2[12]), .CK(clock), .Q(d3[12]) );
  DFF_X1 \d4_reg[12]  ( .D(d3[12]), .CK(clock), .Q(d4[12]) );
  DFF_X1 \d5_reg[12]  ( .D(d4[12]), .CK(clock), .Q(d5[12]) );
  DFF_X1 \d6_reg[12]  ( .D(d5[12]), .CK(clock), .Q(d6[12]) );
  DFF_X1 \d7_reg[12]  ( .D(d6[12]), .CK(clock), .Q(d7[12]) );
  DFF_X1 \d8_reg[12]  ( .D(d7[12]), .CK(clock), .Q(d8[12]) );
  DFF_X1 \d9_reg[12]  ( .D(d8[12]), .CK(clock), .Q(d9[12]) );
  DFF_X1 \d10_reg[12]  ( .D(d9[12]), .CK(clock), .Q(d10[12]) );
  DFF_X1 \d11_reg[12]  ( .D(d10[12]), .CK(clock), .Q(d11[12]) );
  DFF_X1 \d12_reg[12]  ( .D(d11[12]), .CK(clock), .Q(d12[12]) );
  DFF_X1 \d13_reg[12]  ( .D(d12[12]), .CK(clock), .Q(d13[12]) );
  DFF_X1 \d14_reg[12]  ( .D(d13[12]), .CK(clock), .Q(d14[12]) );
  DFF_X1 \d15_reg[12]  ( .D(d14[12]), .CK(clock), .QN(n26) );
  DFF_X1 \d1_reg[11]  ( .D(outA[11]), .CK(clock), .Q(d1[11]) );
  DFF_X1 \d2_reg[11]  ( .D(d1[11]), .CK(clock), .Q(d2[11]) );
  DFF_X1 \d3_reg[11]  ( .D(d2[11]), .CK(clock), .Q(d3[11]) );
  DFF_X1 \d4_reg[11]  ( .D(d3[11]), .CK(clock), .Q(d4[11]) );
  DFF_X1 \d5_reg[11]  ( .D(d4[11]), .CK(clock), .Q(d5[11]) );
  DFF_X1 \d6_reg[11]  ( .D(d5[11]), .CK(clock), .Q(d6[11]) );
  DFF_X1 \d7_reg[11]  ( .D(d6[11]), .CK(clock), .Q(d7[11]) );
  DFF_X1 \d8_reg[11]  ( .D(d7[11]), .CK(clock), .Q(d8[11]) );
  DFF_X1 \d9_reg[11]  ( .D(d8[11]), .CK(clock), .Q(d9[11]) );
  DFF_X1 \d10_reg[11]  ( .D(d9[11]), .CK(clock), .Q(d10[11]) );
  DFF_X1 \d11_reg[11]  ( .D(d10[11]), .CK(clock), .Q(d11[11]) );
  DFF_X1 \d12_reg[11]  ( .D(d11[11]), .CK(clock), .Q(d12[11]) );
  DFF_X1 \d13_reg[11]  ( .D(d12[11]), .CK(clock), .Q(d13[11]) );
  DFF_X1 \d14_reg[11]  ( .D(d13[11]), .CK(clock), .Q(d14[11]) );
  DFF_X1 \d15_reg[11]  ( .D(d14[11]), .CK(clock), .QN(n24) );
  DFF_X1 \d1_reg[10]  ( .D(outA[10]), .CK(clock), .Q(d1[10]) );
  DFF_X1 \d2_reg[10]  ( .D(d1[10]), .CK(clock), .Q(d2[10]) );
  DFF_X1 \d3_reg[10]  ( .D(d2[10]), .CK(clock), .Q(d3[10]) );
  DFF_X1 \d4_reg[10]  ( .D(d3[10]), .CK(clock), .Q(d4[10]) );
  DFF_X1 \d5_reg[10]  ( .D(d4[10]), .CK(clock), .Q(d5[10]) );
  DFF_X1 \d6_reg[10]  ( .D(d5[10]), .CK(clock), .Q(d6[10]) );
  DFF_X1 \d7_reg[10]  ( .D(d6[10]), .CK(clock), .Q(d7[10]) );
  DFF_X1 \d8_reg[10]  ( .D(d7[10]), .CK(clock), .Q(d8[10]) );
  DFF_X1 \d9_reg[10]  ( .D(d8[10]), .CK(clock), .Q(d9[10]) );
  DFF_X1 \d10_reg[10]  ( .D(d9[10]), .CK(clock), .Q(d10[10]) );
  DFF_X1 \d11_reg[10]  ( .D(d10[10]), .CK(clock), .Q(d11[10]) );
  DFF_X1 \d12_reg[10]  ( .D(d11[10]), .CK(clock), .Q(d12[10]) );
  DFF_X1 \d13_reg[10]  ( .D(d12[10]), .CK(clock), .Q(d13[10]) );
  DFF_X1 \d14_reg[10]  ( .D(d13[10]), .CK(clock), .Q(d14[10]) );
  DFF_X1 \d15_reg[10]  ( .D(d14[10]), .CK(clock), .QN(n22) );
  DFF_X1 \d1_reg[9]  ( .D(outA[9]), .CK(clock), .Q(d1[9]) );
  DFF_X1 \d2_reg[9]  ( .D(d1[9]), .CK(clock), .Q(d2[9]) );
  DFF_X1 \d3_reg[9]  ( .D(d2[9]), .CK(clock), .Q(d3[9]) );
  DFF_X1 \d4_reg[9]  ( .D(d3[9]), .CK(clock), .Q(d4[9]) );
  DFF_X1 \d5_reg[9]  ( .D(d4[9]), .CK(clock), .Q(d5[9]) );
  DFF_X1 \d6_reg[9]  ( .D(d5[9]), .CK(clock), .Q(d6[9]) );
  DFF_X1 \d7_reg[9]  ( .D(d6[9]), .CK(clock), .Q(d7[9]) );
  DFF_X1 \d8_reg[9]  ( .D(d7[9]), .CK(clock), .Q(d8[9]) );
  DFF_X1 \d9_reg[9]  ( .D(d8[9]), .CK(clock), .Q(d9[9]) );
  DFF_X1 \d10_reg[9]  ( .D(d9[9]), .CK(clock), .Q(d10[9]) );
  DFF_X1 \d11_reg[9]  ( .D(d10[9]), .CK(clock), .Q(d11[9]) );
  DFF_X1 \d12_reg[9]  ( .D(d11[9]), .CK(clock), .Q(d12[9]) );
  DFF_X1 \d13_reg[9]  ( .D(d12[9]), .CK(clock), .Q(d13[9]) );
  DFF_X1 \d14_reg[9]  ( .D(d13[9]), .CK(clock), .Q(d14[9]) );
  DFF_X1 \d15_reg[9]  ( .D(d14[9]), .CK(clock), .QN(n20) );
  DFF_X1 \d1_reg[8]  ( .D(outA[8]), .CK(clock), .Q(d1[8]) );
  DFF_X1 \d2_reg[8]  ( .D(d1[8]), .CK(clock), .Q(d2[8]) );
  DFF_X1 \d3_reg[8]  ( .D(d2[8]), .CK(clock), .Q(d3[8]) );
  DFF_X1 \d4_reg[8]  ( .D(d3[8]), .CK(clock), .Q(d4[8]) );
  DFF_X1 \d5_reg[8]  ( .D(d4[8]), .CK(clock), .Q(d5[8]) );
  DFF_X1 \d6_reg[8]  ( .D(d5[8]), .CK(clock), .Q(d6[8]) );
  DFF_X1 \d7_reg[8]  ( .D(d6[8]), .CK(clock), .Q(d7[8]) );
  DFF_X1 \d8_reg[8]  ( .D(d7[8]), .CK(clock), .Q(d8[8]) );
  DFF_X1 \d9_reg[8]  ( .D(d8[8]), .CK(clock), .Q(d9[8]) );
  DFF_X1 \d10_reg[8]  ( .D(d9[8]), .CK(clock), .Q(d10[8]) );
  DFF_X1 \d11_reg[8]  ( .D(d10[8]), .CK(clock), .Q(d11[8]) );
  DFF_X1 \d12_reg[8]  ( .D(d11[8]), .CK(clock), .Q(d12[8]) );
  DFF_X1 \d13_reg[8]  ( .D(d12[8]), .CK(clock), .Q(d13[8]) );
  DFF_X1 \d14_reg[8]  ( .D(d13[8]), .CK(clock), .Q(d14[8]) );
  DFF_X1 \d15_reg[8]  ( .D(d14[8]), .CK(clock), .QN(n18) );
  DFF_X1 \d1_reg[7]  ( .D(outA[7]), .CK(clock), .Q(d1[7]) );
  DFF_X1 \d2_reg[7]  ( .D(d1[7]), .CK(clock), .Q(d2[7]) );
  DFF_X1 \d3_reg[7]  ( .D(d2[7]), .CK(clock), .Q(d3[7]) );
  DFF_X1 \d4_reg[7]  ( .D(d3[7]), .CK(clock), .Q(d4[7]) );
  DFF_X1 \d5_reg[7]  ( .D(d4[7]), .CK(clock), .Q(d5[7]) );
  DFF_X1 \d6_reg[7]  ( .D(d5[7]), .CK(clock), .Q(d6[7]) );
  DFF_X1 \d7_reg[7]  ( .D(d6[7]), .CK(clock), .Q(d7[7]) );
  DFF_X1 \d8_reg[7]  ( .D(d7[7]), .CK(clock), .Q(d8[7]) );
  DFF_X1 \d9_reg[7]  ( .D(d8[7]), .CK(clock), .Q(d9[7]) );
  DFF_X1 \d10_reg[7]  ( .D(d9[7]), .CK(clock), .Q(d10[7]) );
  DFF_X1 \d11_reg[7]  ( .D(d10[7]), .CK(clock), .Q(d11[7]) );
  DFF_X1 \d12_reg[7]  ( .D(d11[7]), .CK(clock), .Q(d12[7]) );
  DFF_X1 \d13_reg[7]  ( .D(d12[7]), .CK(clock), .Q(d13[7]) );
  DFF_X1 \d14_reg[7]  ( .D(d13[7]), .CK(clock), .Q(d14[7]) );
  DFF_X1 \d15_reg[7]  ( .D(d14[7]), .CK(clock), .QN(n16) );
  DFF_X1 \d1_reg[6]  ( .D(outA[6]), .CK(clock), .Q(d1[6]) );
  DFF_X1 \d2_reg[6]  ( .D(d1[6]), .CK(clock), .Q(d2[6]) );
  DFF_X1 \d3_reg[6]  ( .D(d2[6]), .CK(clock), .Q(d3[6]) );
  DFF_X1 \d4_reg[6]  ( .D(d3[6]), .CK(clock), .Q(d4[6]) );
  DFF_X1 \d5_reg[6]  ( .D(d4[6]), .CK(clock), .Q(d5[6]) );
  DFF_X1 \d6_reg[6]  ( .D(d5[6]), .CK(clock), .Q(d6[6]) );
  DFF_X1 \d7_reg[6]  ( .D(d6[6]), .CK(clock), .Q(d7[6]) );
  DFF_X1 \d8_reg[6]  ( .D(d7[6]), .CK(clock), .Q(d8[6]) );
  DFF_X1 \d9_reg[6]  ( .D(d8[6]), .CK(clock), .Q(d9[6]) );
  DFF_X1 \d10_reg[6]  ( .D(d9[6]), .CK(clock), .Q(d10[6]) );
  DFF_X1 \d11_reg[6]  ( .D(d10[6]), .CK(clock), .Q(d11[6]) );
  DFF_X1 \d12_reg[6]  ( .D(d11[6]), .CK(clock), .Q(d12[6]) );
  DFF_X1 \d13_reg[6]  ( .D(d12[6]), .CK(clock), .Q(d13[6]) );
  DFF_X1 \d14_reg[6]  ( .D(d13[6]), .CK(clock), .Q(d14[6]) );
  DFF_X1 \d15_reg[6]  ( .D(d14[6]), .CK(clock), .QN(n14) );
  DFF_X1 \d1_reg[5]  ( .D(outA[5]), .CK(clock), .Q(d1[5]) );
  DFF_X1 \d2_reg[5]  ( .D(d1[5]), .CK(clock), .Q(d2[5]) );
  DFF_X1 \d3_reg[5]  ( .D(d2[5]), .CK(clock), .Q(d3[5]) );
  DFF_X1 \d4_reg[5]  ( .D(d3[5]), .CK(clock), .Q(d4[5]) );
  DFF_X1 \d5_reg[5]  ( .D(d4[5]), .CK(clock), .Q(d5[5]) );
  DFF_X1 \d6_reg[5]  ( .D(d5[5]), .CK(clock), .Q(d6[5]) );
  DFF_X1 \d7_reg[5]  ( .D(d6[5]), .CK(clock), .Q(d7[5]) );
  DFF_X1 \d8_reg[5]  ( .D(d7[5]), .CK(clock), .Q(d8[5]) );
  DFF_X1 \d9_reg[5]  ( .D(d8[5]), .CK(clock), .Q(d9[5]) );
  DFF_X1 \d10_reg[5]  ( .D(d9[5]), .CK(clock), .Q(d10[5]) );
  DFF_X1 \d11_reg[5]  ( .D(d10[5]), .CK(clock), .Q(d11[5]) );
  DFF_X1 \d12_reg[5]  ( .D(d11[5]), .CK(clock), .Q(d12[5]) );
  DFF_X1 \d13_reg[5]  ( .D(d12[5]), .CK(clock), .Q(d13[5]) );
  DFF_X1 \d14_reg[5]  ( .D(d13[5]), .CK(clock), .Q(d14[5]) );
  DFF_X1 \d15_reg[5]  ( .D(d14[5]), .CK(clock), .QN(n12) );
  DFF_X1 \d1_reg[4]  ( .D(outA[4]), .CK(clock), .Q(d1[4]) );
  DFF_X1 \d2_reg[4]  ( .D(d1[4]), .CK(clock), .Q(d2[4]) );
  DFF_X1 \d3_reg[4]  ( .D(d2[4]), .CK(clock), .Q(d3[4]) );
  DFF_X1 \d4_reg[4]  ( .D(d3[4]), .CK(clock), .Q(d4[4]) );
  DFF_X1 \d5_reg[4]  ( .D(d4[4]), .CK(clock), .Q(d5[4]) );
  DFF_X1 \d6_reg[4]  ( .D(d5[4]), .CK(clock), .Q(d6[4]) );
  DFF_X1 \d7_reg[4]  ( .D(d6[4]), .CK(clock), .Q(d7[4]) );
  DFF_X1 \d8_reg[4]  ( .D(d7[4]), .CK(clock), .Q(d8[4]) );
  DFF_X1 \d9_reg[4]  ( .D(d8[4]), .CK(clock), .Q(d9[4]) );
  DFF_X1 \d10_reg[4]  ( .D(d9[4]), .CK(clock), .Q(d10[4]) );
  DFF_X1 \d11_reg[4]  ( .D(d10[4]), .CK(clock), .Q(d11[4]) );
  DFF_X1 \d12_reg[4]  ( .D(d11[4]), .CK(clock), .Q(d12[4]) );
  DFF_X1 \d13_reg[4]  ( .D(d12[4]), .CK(clock), .Q(d13[4]) );
  DFF_X1 \d14_reg[4]  ( .D(d13[4]), .CK(clock), .Q(d14[4]) );
  DFF_X1 \d15_reg[4]  ( .D(d14[4]), .CK(clock), .QN(n10) );
  DFF_X1 \d1_reg[3]  ( .D(outA[3]), .CK(clock), .Q(d1[3]) );
  DFF_X1 \d2_reg[3]  ( .D(d1[3]), .CK(clock), .Q(d2[3]) );
  DFF_X1 \d3_reg[3]  ( .D(d2[3]), .CK(clock), .Q(d3[3]) );
  DFF_X1 \d4_reg[3]  ( .D(d3[3]), .CK(clock), .Q(d4[3]) );
  DFF_X1 \d5_reg[3]  ( .D(d4[3]), .CK(clock), .Q(d5[3]) );
  DFF_X1 \d6_reg[3]  ( .D(d5[3]), .CK(clock), .Q(d6[3]) );
  DFF_X1 \d7_reg[3]  ( .D(d6[3]), .CK(clock), .Q(d7[3]) );
  DFF_X1 \d8_reg[3]  ( .D(d7[3]), .CK(clock), .Q(d8[3]) );
  DFF_X1 \d9_reg[3]  ( .D(d8[3]), .CK(clock), .Q(d9[3]) );
  DFF_X1 \d10_reg[3]  ( .D(d9[3]), .CK(clock), .Q(d10[3]) );
  DFF_X1 \d11_reg[3]  ( .D(d10[3]), .CK(clock), .Q(d11[3]) );
  DFF_X1 \d12_reg[3]  ( .D(d11[3]), .CK(clock), .Q(d12[3]) );
  DFF_X1 \d13_reg[3]  ( .D(d12[3]), .CK(clock), .Q(d13[3]) );
  DFF_X1 \d14_reg[3]  ( .D(d13[3]), .CK(clock), .Q(d14[3]) );
  DFF_X1 \d15_reg[3]  ( .D(d14[3]), .CK(clock), .QN(n8) );
  DFF_X1 \d1_reg[2]  ( .D(outA[2]), .CK(clock), .Q(d1[2]) );
  DFF_X1 \d2_reg[2]  ( .D(d1[2]), .CK(clock), .Q(d2[2]) );
  DFF_X1 \d3_reg[2]  ( .D(d2[2]), .CK(clock), .Q(d3[2]) );
  DFF_X1 \d4_reg[2]  ( .D(d3[2]), .CK(clock), .Q(d4[2]) );
  DFF_X1 \d5_reg[2]  ( .D(d4[2]), .CK(clock), .Q(d5[2]) );
  DFF_X1 \d6_reg[2]  ( .D(d5[2]), .CK(clock), .Q(d6[2]) );
  DFF_X1 \d7_reg[2]  ( .D(d6[2]), .CK(clock), .Q(d7[2]) );
  DFF_X1 \d8_reg[2]  ( .D(d7[2]), .CK(clock), .Q(d8[2]) );
  DFF_X1 \d9_reg[2]  ( .D(d8[2]), .CK(clock), .Q(d9[2]) );
  DFF_X1 \d10_reg[2]  ( .D(d9[2]), .CK(clock), .Q(d10[2]) );
  DFF_X1 \d11_reg[2]  ( .D(d10[2]), .CK(clock), .Q(d11[2]) );
  DFF_X1 \d12_reg[2]  ( .D(d11[2]), .CK(clock), .Q(d12[2]) );
  DFF_X1 \d13_reg[2]  ( .D(d12[2]), .CK(clock), .Q(d13[2]) );
  DFF_X1 \d14_reg[2]  ( .D(d13[2]), .CK(clock), .Q(d14[2]) );
  DFF_X1 \d15_reg[2]  ( .D(d14[2]), .CK(clock), .QN(n6) );
  DFF_X1 \d1_reg[1]  ( .D(outA[1]), .CK(clock), .Q(d1[1]) );
  DFF_X1 \d2_reg[1]  ( .D(d1[1]), .CK(clock), .Q(d2[1]) );
  DFF_X1 \d3_reg[1]  ( .D(d2[1]), .CK(clock), .Q(d3[1]) );
  DFF_X1 \d4_reg[1]  ( .D(d3[1]), .CK(clock), .Q(d4[1]) );
  DFF_X1 \d5_reg[1]  ( .D(d4[1]), .CK(clock), .Q(d5[1]) );
  DFF_X1 \d6_reg[1]  ( .D(d5[1]), .CK(clock), .Q(d6[1]) );
  DFF_X1 \d7_reg[1]  ( .D(d6[1]), .CK(clock), .Q(d7[1]) );
  DFF_X1 \d8_reg[1]  ( .D(d7[1]), .CK(clock), .Q(d8[1]) );
  DFF_X1 \d9_reg[1]  ( .D(d8[1]), .CK(clock), .Q(d9[1]) );
  DFF_X1 \d10_reg[1]  ( .D(d9[1]), .CK(clock), .Q(d10[1]) );
  DFF_X1 \d11_reg[1]  ( .D(d10[1]), .CK(clock), .Q(d11[1]) );
  DFF_X1 \d12_reg[1]  ( .D(d11[1]), .CK(clock), .Q(d12[1]) );
  DFF_X1 \d13_reg[1]  ( .D(d12[1]), .CK(clock), .Q(d13[1]) );
  DFF_X1 \d14_reg[1]  ( .D(d13[1]), .CK(clock), .Q(d14[1]) );
  DFF_X1 \d15_reg[1]  ( .D(d14[1]), .CK(clock), .QN(n4) );
  DFF_X1 \d1_reg[0]  ( .D(outA[0]), .CK(clock), .Q(d1[0]) );
  DFF_X1 \d2_reg[0]  ( .D(d1[0]), .CK(clock), .Q(d2[0]) );
  DFF_X1 \d3_reg[0]  ( .D(d2[0]), .CK(clock), .Q(d3[0]) );
  DFF_X1 \d4_reg[0]  ( .D(d3[0]), .CK(clock), .Q(d4[0]) );
  DFF_X1 \d5_reg[0]  ( .D(d4[0]), .CK(clock), .Q(d5[0]) );
  DFF_X1 \d6_reg[0]  ( .D(d5[0]), .CK(clock), .Q(d6[0]) );
  DFF_X1 \d7_reg[0]  ( .D(d6[0]), .CK(clock), .Q(d7[0]) );
  DFF_X1 \d8_reg[0]  ( .D(d7[0]), .CK(clock), .Q(d8[0]) );
  DFF_X1 \d9_reg[0]  ( .D(d8[0]), .CK(clock), .Q(d9[0]) );
  DFF_X1 \d10_reg[0]  ( .D(d9[0]), .CK(clock), .Q(d10[0]) );
  DFF_X1 \d11_reg[0]  ( .D(d10[0]), .CK(clock), .Q(d11[0]) );
  DFF_X1 \d12_reg[0]  ( .D(d11[0]), .CK(clock), .Q(d12[0]) );
  DFF_X1 \d13_reg[0]  ( .D(d12[0]), .CK(clock), .Q(d13[0]) );
  DFF_X1 \d14_reg[0]  ( .D(d13[0]), .CK(clock), .Q(d14[0]) );
  DFF_X1 \d15_reg[0]  ( .D(d14[0]), .CK(clock), .QN(n2) );
  OAI22_X2 U3 ( .A1(n2), .A2(n903), .B1(n3), .B2(n902), .ZN(n98) );
  OAI22_X2 U4 ( .A1(n4), .A2(n903), .B1(n5), .B2(n902), .ZN(n99) );
  OAI22_X2 U5 ( .A1(n6), .A2(n903), .B1(n7), .B2(adder_output[24]), .ZN(n100)
         );
  OAI22_X2 U6 ( .A1(n8), .A2(n903), .B1(n9), .B2(n902), .ZN(n101) );
  OAI22_X2 U7 ( .A1(n10), .A2(n903), .B1(n11), .B2(n902), .ZN(n102) );
  OAI22_X2 U8 ( .A1(n12), .A2(n903), .B1(n13), .B2(adder_output[24]), .ZN(n103) );
  OAI22_X2 U9 ( .A1(n14), .A2(n903), .B1(n15), .B2(n902), .ZN(n104) );
  OAI22_X2 U10 ( .A1(n16), .A2(n903), .B1(n17), .B2(n902), .ZN(n105) );
  OAI22_X2 U11 ( .A1(n18), .A2(n903), .B1(n19), .B2(adder_output[24]), .ZN(
        n106) );
  OAI22_X2 U12 ( .A1(n20), .A2(n903), .B1(n21), .B2(n902), .ZN(n107) );
  OAI22_X2 U13 ( .A1(n22), .A2(n903), .B1(n23), .B2(n902), .ZN(n108) );
  OAI22_X2 U14 ( .A1(n24), .A2(n903), .B1(n25), .B2(adder_output[24]), .ZN(
        n109) );
  OAI22_X2 U15 ( .A1(n26), .A2(n903), .B1(n27), .B2(n902), .ZN(n110) );
  OAI22_X2 U16 ( .A1(n28), .A2(n903), .B1(n29), .B2(n902), .ZN(n111) );
  OAI22_X2 U17 ( .A1(n30), .A2(n903), .B1(n31), .B2(n902), .ZN(n112) );
  OAI22_X2 U18 ( .A1(n32), .A2(n903), .B1(n33), .B2(adder_output[24]), .ZN(
        n113) );
  OAI22_X2 U19 ( .A1(n34), .A2(n903), .B1(n35), .B2(n902), .ZN(n114) );
  OAI22_X2 U20 ( .A1(n36), .A2(n903), .B1(n37), .B2(adder_output[24]), .ZN(
        n115) );
  OAI22_X2 U21 ( .A1(n38), .A2(n903), .B1(n39), .B2(n902), .ZN(n116) );
  OAI22_X2 U22 ( .A1(n40), .A2(n903), .B1(n41), .B2(adder_output[24]), .ZN(
        n117) );
  OAI22_X2 U23 ( .A1(n42), .A2(n903), .B1(n43), .B2(n902), .ZN(n118) );
  OAI22_X2 U24 ( .A1(n44), .A2(n903), .B1(n45), .B2(adder_output[24]), .ZN(
        n119) );
  OAI22_X2 U25 ( .A1(n46), .A2(n903), .B1(n47), .B2(n902), .ZN(n120) );
  OAI22_X2 U26 ( .A1(n48), .A2(n903), .B1(n49), .B2(adder_output[24]), .ZN(
        n121) );
  OAI22_X2 U27 ( .A1(n50), .A2(n903), .B1(n51), .B2(n902), .ZN(n122) );
  OAI22_X2 U28 ( .A1(n52), .A2(n903), .B1(n53), .B2(n902), .ZN(n123) );
  OAI22_X2 U29 ( .A1(n54), .A2(n903), .B1(n55), .B2(n902), .ZN(n124) );
  OAI22_X2 U30 ( .A1(n56), .A2(n903), .B1(n57), .B2(n902), .ZN(n125) );
  OAI22_X2 U31 ( .A1(n58), .A2(n903), .B1(n59), .B2(n902), .ZN(n126) );
  OAI22_X2 U32 ( .A1(n60), .A2(n903), .B1(n61), .B2(n902), .ZN(n127) );
  OAI22_X2 U33 ( .A1(n62), .A2(n903), .B1(n63), .B2(n902), .ZN(n128) );
  OAI22_X2 U34 ( .A1(n64), .A2(n903), .B1(n65), .B2(n902), .ZN(n129) );
  OAI22_X2 U35 ( .A1(n66), .A2(n903), .B1(n67), .B2(n902), .ZN(n130) );
  OAI22_X2 U36 ( .A1(n68), .A2(n903), .B1(n69), .B2(n902), .ZN(n131) );
  OAI22_X2 U37 ( .A1(n70), .A2(n903), .B1(n71), .B2(n902), .ZN(n132) );
  OAI22_X2 U38 ( .A1(n72), .A2(n903), .B1(n73), .B2(n902), .ZN(n133) );
  OAI22_X2 U39 ( .A1(n74), .A2(n903), .B1(n75), .B2(adder_output[24]), .ZN(
        n134) );
  OAI22_X2 U40 ( .A1(n76), .A2(n903), .B1(n77), .B2(adder_output[24]), .ZN(
        n135) );
  OAI22_X2 U41 ( .A1(n78), .A2(n903), .B1(n79), .B2(n902), .ZN(n136) );
  OAI22_X2 U42 ( .A1(n80), .A2(n903), .B1(n81), .B2(n902), .ZN(n137) );
  OAI22_X2 U43 ( .A1(n82), .A2(n903), .B1(n83), .B2(n902), .ZN(n138) );
  OAI22_X2 U44 ( .A1(n84), .A2(n903), .B1(n85), .B2(n902), .ZN(n139) );
  OAI22_X2 U45 ( .A1(n86), .A2(n903), .B1(n87), .B2(n902), .ZN(n140) );
  OAI22_X2 U46 ( .A1(n88), .A2(n903), .B1(n89), .B2(n902), .ZN(n141) );
  OAI22_X2 U47 ( .A1(n90), .A2(n903), .B1(n91), .B2(n902), .ZN(n142) );
  OAI22_X2 U48 ( .A1(n92), .A2(n903), .B1(n93), .B2(n902), .ZN(n143) );
  OAI22_X2 U49 ( .A1(n94), .A2(n903), .B1(n95), .B2(n902), .ZN(n144) );
  OAI22_X2 U50 ( .A1(n96), .A2(n903), .B1(n97), .B2(n902), .ZN(n145) );
  update_1 u2 ( .X({X[15:8], n803, n801, n799, n797, n795, n793, n791, n789}), 
        .Y({Y[15:8], n787, n785, n783, n781, n779, n777, n775, n773}), 
        .Y_ramX(Y_ramX), .Y_ramY(Y_ramY) );
  update_2 u4 ( .X({X[15:8], n803, n801, n799, n797, n795, n793, n791, n789}), 
        .Y({Y[15:8], n787, n785, n783, n781, n779, n777, n775, n773}), .RowX(
        RowX), .RowY(RowY), .Y_ramX(Y_ramX), .Y_ramY(Y_ramY), .Row_noX(Row_noX), .Row_noY(Row_noY), .clock(clock), .EnableChange(EnableChange), .FoundX(
        FoundX), .FoundY(FoundY), .FlagX(FlagX), .FlagY(FlagY), 
        .DiagonalDoneX(DiagonalDoneX), .DiagonalDoneY(DiagonalDoneY), .WireX(
        WireX), .WireY(WireY) );
  MainArbiter_1 u15 ( .reset(n901), .clock(clock), .EnableChange(EnableChange), 
        .Update_1Req1(Y_ramX), .Update_1Req2(Y_ramY), .Update_2Req1(Row_noX), 
        .Update_2Req2(Row_noY), .Row1({n771, n769, n767, n765, n763, n761, 
        n759, n757, n755, n753, n751, n749, n747, n745, n743, n741, 
        ReadBus1[239:192], n739, n737, n735, n733, n731, n729, n727, n725, 
        n723, n721, n719, n717, n715, n713, n711, n709, ReadBus1[175:128], 
        n707, n705, n703, n701, n699, n697, n695, n693, n691, n689, n687, n685, 
        n683, n681, n679, n677, ReadBus1[111:107], n675, n673, n671, n669, 
        n667, n665, n663, n661, n659, n657, n655, ReadBus1[95:91], n653, n651, 
        n649, n647, n645, n643, n641, n639, n637, n635, n633, ReadBus1[79:75], 
        n631, n629, n627, n625, n623, n621, n619, n617, n615, n613, n611, n609, 
        n607, n605, n603, n601, n599, n597, n595, n593, n591, n589, n587, n585, 
        n583, n581, n579, ReadBus1[47:0]}), .Row2(ReadBus2), .OutputReq1(
        ReadAddress1), .OutputReq2(ReadAddress2), .Output_1Row1(RowX), 
        .Output_1Row2(RowY), .Output_2Row1(NewRowX), .Output_2Row2(NewRowY), 
        .FlagX(FlagX), .FlagY(FlagY), .DiagonalDoneX(DiagonalXDone), 
        .DiagonalDoneY(1'b1), .WE(WE), .PosDX(PosDX), .PaddedRow(PaddedRow), 
        .WriteReq(WriteReq), .WriteBus(WriteBus), .NewDiagonalX(NewDiagonalX), 
        .NewDiagonalY(NewDiagonalY), .NewElement(NewElement), .ArbiterElement(
        ArbiterElement), .ArbiterPos(ArbiterPos), .OutputPaddedRow(
        OutputPaddedRow), .PosDY(PosDY), .PosRowX(PosRowX), .PosRowY(PosRowY), 
        .ComputeReq(ComputeReq), .OutputCompute(OutputCompute), .CompStart(
        CompStart), .EOC_Flag(EOC_Flag) );
  update_3 u6 ( .reset(n901), .clock(clock), .X({X[15:8], n803, n801, n799, 
        n797, n795, n793, n791, n789}), .Y({Y[15:8], n787, n785, n783, n781, 
        n779, n777, n775, n773}), .NewRowX(NewRowX), .NewRowY(NewRowY), 
        .DiagonalX(DiagonalX), .DiagonalY(DiagonalY), .PosDX(PosDX), .PosDY(
        PosDY), .DiagonalDoneX(DiagonalDoneX), .DiagonalDoneY(DiagonalDoneY), 
        .Row_noX(Row_noX), .Row_noY(Row_noY), .EnableChange(EnableChange) );
  update_3_1 u7 ( .reset(n901), .clock(clock), .X({X[15:8], n803, n801, n799, 
        n797, n795, n793, n791, n789}), .Y({Y[15:8], n787, n785, n783, n781, 
        n779, n777, n775, n773}), .NewRowX(NewRowX), .NewRowY(NewRowY), 
        .Element(ElementUpdate), .PosRowX(PosRowX), .PosRowY(PosRowY), .PosDX(
        PosDX), .PosDY(PosDY), .FoundX(FoundX), .FoundY(FoundY), .Row_noX(
        Row_noX), .Row_noY(Row_noY), .DiagonalDoneX(DiagonalDoneX), 
        .DiagonalDoneY(DiagonalDoneY), .EnableChange(EnableChange), .WireX(
        WireX), .WireY(WireY) );
  arithController u8 ( .clock(clock), .reset(n901), .DiagonalX(DiagonalX), 
        .DiagonalY(DiagonalY), .Element(ElementUpdate), .NewElement(NewElement), .EnableChange(EnableChange), .SubInput1(SubInput1), .SubInput2(SubInput2), 
        .AddInput1(AddInput1), .AddInput2(AddInput2), .NewDiagonalX(
        NewDiagonalX), .NewDiagonalY(NewDiagonalY), .SubOutput(SubOutput), 
        .AddOutput(AddOutput), .DiagonalXDone(DiagonalXDone) );
  pad_3 u11 ( .Element(ArbiterElement), .PosElement(ArbiterPos), .Y_ramRow(
        OutputPaddedRow), .PaddedRow(PaddedRow) );
  selector a1 ( .dataY(OutputCompute), .count({SYNOPSYS_UNCONNECTED__0, 
        count[1:0]}), .EOF(EOF) );
  EOF_reg a31 ( .clock(clock), .reset(n901), .EOF(EOF), .sig(sig_OP) );
  y_arbiter a2 ( .reset(n901), .clock(clock), .addressY(ComputeReq), .count2({
        1'b0, count[1:0]}), .EOF(EOF), .MainCount({SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, \MainCount1[0] }), .sig(sig_OP), .EOC_Flag(
        EOC_Flag), .CompStart(CompStart) );
  decoder a3 ( .clock(clock), .reset(n901), .data(OutputCompute), .Diagonal(
        outA), .Element(outB), .ElementAddr(ElementAddr), .EOF(EOF), .sig(
        sig_OP), .CompStart(CompStart) );
  v_arbiter a5 ( .vop1(vop1), .vop2(vop2), .vop3(vop3), .vop4(vop4), .rowno(
        ElementAddr), .clock(clock), .Vout(Vout), .Rowread1(Rowread1), 
        .Rowread2(Rowread2), .Rowread3(Rowread3), .Rowread4(Rowread4), 
        .count2(\MainCount1[0] ) );
  sync a10 ( .clock(clock), .ElementY(outB), .ElementV(Vout), .SyncY(SyncY), 
        .SyncV(SyncV) );
  syncDiv a9 ( .element1(diagOut), .op1(diagonalC), .op2(diagonalD), .clock(
        clock) );
  syncMult a4 ( .clock(clock), .SyncY(SyncY), .SyncMultY(SyncMultY), 
        .multinput({n899, n897, n895, n893, n891, n889, n887, n885, n883, n881, 
        n879, n877, n875, n873, n871, n869, n867, n865, n863, n861, n859, n857, 
        n855, n853, n851, n849, n847, n845, n843, n841, n839, n837, n835, n833, 
        n831, n829, n827, n825, n823, n821, n819, n817, n815, n813, n811, n809, 
        n807, n805}), .mult_output(mult_output) );
  controller2_1 a12 ( .clock(clock), .reset(n901), .accum_in({n902, 
        adder_output[23:0]}), .feedback(adder_input), .set_bit(mult_output[48]), .element(mult_output[48:24]) );
  syncAccum_0 a14 ( .clock(clock), .mult_output(mult_output[48:24]), 
        .accum_input(accum_input), .accum_output(accum_output), 
        .accum_output25(adder_output) );
  controller2_0 a26 ( .clock(clock), .reset(n901), .accum_in(adder_output_imag), .feedback(adder_input_imag), .set_bit(mult_output[48]), .element({
        mult_output[48], mult_output[23:0]}) );
  syncAccum_1 a15 ( .clock(clock), .mult_output({mult_output[48], 
        mult_output[23:0]}), .accum_input(accum_input_imag), .accum_output(
        accum_output_imag), .accum_output25(adder_output_imag) );
  isched a17 ( .clock(clock), .reset(n901), .addressI(addressI), .data(outI), 
        .dataI(dataI), .FinalOutput(adder_out7), .sig(sig_OP) );
  write_enable a24 ( .input_data(op_final), .input_data2(op_reg), .signal(
        signal), .signal2(signal2) );
  v_sched a25 ( .signal(signal), .signal2(signal2), .clock(clock), .reset(n901), .write_addr1(write_addr1), .we1(we1), .write_addr2(write_addr2), .we2(we2), 
        .write_addr3(write_addr3), .we3(we3), .write_addr4(write_addr4), .we4(
        we4), .sig_I(sig_OP), .count2(\MainCount1[0] ) );
  DFF_X2 \op_reg_reg[14]  ( .D(op_final[14]), .CK(clock), .Q(op_reg[14]) );
  DFF_X2 \op_reg_reg[17]  ( .D(op_final[17]), .CK(clock), .Q(op_reg[17]) );
  DFF_X2 \op_reg_reg[4]  ( .D(op_final[4]), .CK(clock), .Q(op_reg[4]) );
  DFF_X2 \op_reg_reg[7]  ( .D(op_final[7]), .CK(clock), .Q(op_reg[7]) );
  DFF_X2 \op_reg_reg[22]  ( .D(op_final[22]), .CK(clock), .Q(op_reg[22]) );
  DFF_X2 \op_reg_reg[25]  ( .D(op_final[25]), .CK(clock), .Q(op_reg[25]) );
  DFF_X2 \op_reg_reg[28]  ( .D(op_final[28]), .CK(clock), .Q(op_reg[28]) );
  DFF_X2 \op_reg_reg[33]  ( .D(op_final[33]), .CK(clock), .Q(op_reg[33]) );
  DFF_X2 \op_reg_reg[36]  ( .D(op_final[36]), .CK(clock), .Q(op_reg[36]) );
  DFF_X2 \op_reg_reg[39]  ( .D(op_final[39]), .CK(clock), .Q(op_reg[39]) );
  DFF_X2 \op_reg_reg[44]  ( .D(op_final[44]), .CK(clock), .Q(op_reg[44]) );
  DFF_X2 \op_reg_reg[1]  ( .D(op_final[1]), .CK(clock), .Q(op_reg[1]) );
  DFF_X2 \op_reg_reg[11]  ( .D(op_final[11]), .CK(clock), .Q(op_reg[11]) );
  DFF_X2 \op_reg_reg[30]  ( .D(op_final[30]), .CK(clock), .Q(op_reg[30]) );
  DFF_X2 \op_reg_reg[41]  ( .D(op_final[41]), .CK(clock), .Q(op_reg[41]) );
  DFF_X2 \op_reg_reg[15]  ( .D(op_final[15]), .CK(clock), .Q(op_reg[15]) );
  DFF_X2 \op_reg_reg[3]  ( .D(op_final[3]), .CK(clock), .Q(op_reg[3]) );
  DFF_X2 \op_reg_reg[5]  ( .D(op_final[5]), .CK(clock), .Q(op_reg[5]) );
  DFF_X2 \op_reg_reg[23]  ( .D(op_final[23]), .CK(clock), .Q(op_reg[23]) );
  DFF_X2 \op_reg_reg[12]  ( .D(op_final[12]), .CK(clock), .Q(op_reg[12]) );
  DFF_X2 \op_reg_reg[20]  ( .D(op_final[20]), .CK(clock), .Q(op_reg[20]) );
  DFF_X2 \op_reg_reg[31]  ( .D(op_final[31]), .CK(clock), .Q(op_reg[31]) );
  DFF_X2 \op_reg_reg[42]  ( .D(op_final[42]), .CK(clock), .Q(op_reg[42]) );
  DFF_X2 \diagOut_reg[0]  ( .D(n98), .CK(clock), .Q(diagOut[0]), .QN(n3) );
  DFF_X2 \diagOut_reg[1]  ( .D(n99), .CK(clock), .Q(diagOut[1]), .QN(n5) );
  DFF_X2 \diagOut_reg[2]  ( .D(n100), .CK(clock), .Q(diagOut[2]), .QN(n7) );
  DFF_X2 \diagOut_reg[3]  ( .D(n101), .CK(clock), .Q(diagOut[3]), .QN(n9) );
  DFF_X2 \diagOut_reg[4]  ( .D(n102), .CK(clock), .Q(diagOut[4]), .QN(n11) );
  DFF_X2 \diagOut_reg[5]  ( .D(n103), .CK(clock), .Q(diagOut[5]), .QN(n13) );
  DFF_X2 \diagOut_reg[6]  ( .D(n104), .CK(clock), .Q(diagOut[6]), .QN(n15) );
  DFF_X2 \diagOut_reg[7]  ( .D(n105), .CK(clock), .Q(diagOut[7]), .QN(n17) );
  DFF_X2 \diagOut_reg[8]  ( .D(n106), .CK(clock), .Q(diagOut[8]), .QN(n19) );
  DFF_X2 \diagOut_reg[9]  ( .D(n107), .CK(clock), .Q(diagOut[9]), .QN(n21) );
  DFF_X2 \diagOut_reg[10]  ( .D(n108), .CK(clock), .Q(diagOut[10]), .QN(n23)
         );
  DFF_X2 \diagOut_reg[11]  ( .D(n109), .CK(clock), .Q(diagOut[11]), .QN(n25)
         );
  DFF_X2 \diagOut_reg[12]  ( .D(n110), .CK(clock), .Q(diagOut[12]), .QN(n27)
         );
  DFF_X2 \diagOut_reg[13]  ( .D(n111), .CK(clock), .Q(diagOut[13]), .QN(n29)
         );
  DFF_X2 \diagOut_reg[14]  ( .D(n112), .CK(clock), .Q(diagOut[14]), .QN(n31)
         );
  DFF_X2 \diagOut_reg[15]  ( .D(n113), .CK(clock), .Q(diagOut[15]), .QN(n33)
         );
  DFF_X2 \diagOut_reg[16]  ( .D(n114), .CK(clock), .Q(diagOut[16]), .QN(n35)
         );
  DFF_X2 \diagOut_reg[17]  ( .D(n115), .CK(clock), .Q(diagOut[17]), .QN(n37)
         );
  DFF_X2 \diagOut_reg[18]  ( .D(n116), .CK(clock), .Q(diagOut[18]), .QN(n39)
         );
  DFF_X2 \diagOut_reg[19]  ( .D(n117), .CK(clock), .Q(diagOut[19]), .QN(n41)
         );
  DFF_X2 \diagOut_reg[20]  ( .D(n118), .CK(clock), .Q(diagOut[20]), .QN(n43)
         );
  DFF_X2 \diagOut_reg[21]  ( .D(n119), .CK(clock), .Q(diagOut[21]), .QN(n45)
         );
  DFF_X2 \diagOut_reg[22]  ( .D(n120), .CK(clock), .Q(diagOut[22]), .QN(n47)
         );
  DFF_X2 \diagOut_reg[23]  ( .D(n121), .CK(clock), .Q(diagOut[23]), .QN(n49)
         );
  DFF_X2 \diagOut_reg[24]  ( .D(n122), .CK(clock), .Q(diagOut[24]), .QN(n51)
         );
  DFF_X2 \diagOut_reg[25]  ( .D(n123), .CK(clock), .Q(diagOut[25]), .QN(n53)
         );
  DFF_X2 \diagOut_reg[26]  ( .D(n124), .CK(clock), .Q(diagOut[26]), .QN(n55)
         );
  DFF_X2 \diagOut_reg[27]  ( .D(n125), .CK(clock), .Q(diagOut[27]), .QN(n57)
         );
  DFF_X2 \diagOut_reg[28]  ( .D(n126), .CK(clock), .Q(diagOut[28]), .QN(n59)
         );
  DFF_X2 \diagOut_reg[29]  ( .D(n127), .CK(clock), .Q(diagOut[29]), .QN(n61)
         );
  DFF_X2 \diagOut_reg[30]  ( .D(n128), .CK(clock), .Q(diagOut[30]), .QN(n63)
         );
  DFF_X2 \diagOut_reg[31]  ( .D(n129), .CK(clock), .Q(diagOut[31]), .QN(n65)
         );
  DFF_X2 \diagOut_reg[32]  ( .D(n130), .CK(clock), .Q(diagOut[32]), .QN(n67)
         );
  DFF_X2 \diagOut_reg[33]  ( .D(n131), .CK(clock), .Q(diagOut[33]), .QN(n69)
         );
  DFF_X2 \diagOut_reg[34]  ( .D(n132), .CK(clock), .Q(diagOut[34]), .QN(n71)
         );
  DFF_X2 \diagOut_reg[35]  ( .D(n133), .CK(clock), .Q(diagOut[35]), .QN(n73)
         );
  DFF_X2 \diagOut_reg[36]  ( .D(n134), .CK(clock), .Q(diagOut[36]), .QN(n75)
         );
  DFF_X2 \diagOut_reg[37]  ( .D(n135), .CK(clock), .Q(diagOut[37]), .QN(n77)
         );
  DFF_X2 \diagOut_reg[38]  ( .D(n136), .CK(clock), .Q(diagOut[38]), .QN(n79)
         );
  DFF_X2 \diagOut_reg[39]  ( .D(n137), .CK(clock), .Q(diagOut[39]), .QN(n81)
         );
  DFF_X2 \diagOut_reg[40]  ( .D(n138), .CK(clock), .Q(diagOut[40]), .QN(n83)
         );
  DFF_X2 \diagOut_reg[41]  ( .D(n139), .CK(clock), .Q(diagOut[41]), .QN(n85)
         );
  DFF_X2 \diagOut_reg[42]  ( .D(n140), .CK(clock), .Q(diagOut[42]), .QN(n87)
         );
  DFF_X2 \diagOut_reg[43]  ( .D(n141), .CK(clock), .Q(diagOut[43]), .QN(n89)
         );
  DFF_X2 \diagOut_reg[44]  ( .D(n142), .CK(clock), .Q(diagOut[44]), .QN(n91)
         );
  DFF_X2 \diagOut_reg[45]  ( .D(n143), .CK(clock), .Q(diagOut[45]), .QN(n93)
         );
  DFF_X2 \diagOut_reg[46]  ( .D(n144), .CK(clock), .Q(diagOut[46]), .QN(n95)
         );
  DFF_X2 \diagOut_reg[47]  ( .D(n145), .CK(clock), .Q(diagOut[47]), .QN(n97)
         );
  DFF_X2 \op_reg_reg[47]  ( .D(op_final[47]), .CK(clock), .Q(op_reg[47]) );
  DFF_X2 \delay1_reg[0]  ( .D(adder_out7_imag[0]), .CK(clock), .Q(delay1[0])
         );
  DFF_X2 \delay1_reg[1]  ( .D(adder_out7_imag[1]), .CK(clock), .Q(delay1[1])
         );
  DFF_X2 \delay1_reg[2]  ( .D(adder_out7_imag[2]), .CK(clock), .Q(delay1[2])
         );
  DFF_X2 \delay1_reg[3]  ( .D(adder_out7_imag[3]), .CK(clock), .Q(delay1[3])
         );
  DFF_X2 \delay1_reg[4]  ( .D(adder_out7_imag[4]), .CK(clock), .Q(delay1[4])
         );
  DFF_X2 \delay1_reg[5]  ( .D(adder_out7_imag[5]), .CK(clock), .Q(delay1[5])
         );
  DFF_X2 \delay1_reg[6]  ( .D(adder_out7_imag[6]), .CK(clock), .Q(delay1[6])
         );
  DFF_X2 \delay1_reg[7]  ( .D(adder_out7_imag[7]), .CK(clock), .Q(delay1[7])
         );
  DFF_X2 \delay1_reg[8]  ( .D(adder_out7_imag[8]), .CK(clock), .Q(delay1[8])
         );
  DFF_X2 \delay1_reg[9]  ( .D(adder_out7_imag[9]), .CK(clock), .Q(delay1[9])
         );
  DFF_X2 \delay1_reg[10]  ( .D(adder_out7_imag[10]), .CK(clock), .Q(delay1[10]) );
  DFF_X2 \delay1_reg[11]  ( .D(adder_out7_imag[11]), .CK(clock), .Q(delay1[11]) );
  DFF_X2 \delay1_reg[12]  ( .D(adder_out7_imag[12]), .CK(clock), .Q(delay1[12]) );
  DFF_X2 \delay1_reg[13]  ( .D(adder_out7_imag[13]), .CK(clock), .Q(delay1[13]) );
  DFF_X2 \delay1_reg[14]  ( .D(adder_out7_imag[14]), .CK(clock), .Q(delay1[14]) );
  DFF_X2 \delay1_reg[15]  ( .D(adder_out7_imag[15]), .CK(clock), .Q(delay1[15]) );
  DFF_X2 \delay1_reg[16]  ( .D(adder_out7_imag[16]), .CK(clock), .Q(delay1[16]) );
  DFF_X2 \delay1_reg[17]  ( .D(adder_out7_imag[17]), .CK(clock), .Q(delay1[17]) );
  DFF_X2 \delay1_reg[18]  ( .D(adder_out7_imag[18]), .CK(clock), .Q(delay1[18]) );
  DFF_X2 \delay1_reg[19]  ( .D(adder_out7_imag[19]), .CK(clock), .Q(delay1[19]) );
  DFF_X2 \delay1_reg[20]  ( .D(adder_out7_imag[20]), .CK(clock), .Q(delay1[20]) );
  DFF_X2 \delay1_reg[21]  ( .D(adder_out7_imag[21]), .CK(clock), .Q(delay1[21]) );
  DFF_X2 \delay1_reg[22]  ( .D(adder_out7_imag[22]), .CK(clock), .Q(delay1[22]) );
  DFF_X2 \delay1_reg[23]  ( .D(adder_out7_imag[23]), .CK(clock), .Q(delay1[23]) );
  DFF_X2 \delay1_reg[24]  ( .D(adder_out7[0]), .CK(clock), .Q(delay1[24]) );
  DFF_X2 \delay1_reg[25]  ( .D(adder_out7[1]), .CK(clock), .Q(delay1[25]) );
  DFF_X2 \delay1_reg[26]  ( .D(adder_out7[2]), .CK(clock), .Q(delay1[26]) );
  DFF_X2 \delay1_reg[27]  ( .D(adder_out7[3]), .CK(clock), .Q(delay1[27]) );
  DFF_X2 \delay1_reg[28]  ( .D(adder_out7[4]), .CK(clock), .Q(delay1[28]) );
  DFF_X2 \delay1_reg[29]  ( .D(adder_out7[5]), .CK(clock), .Q(delay1[29]) );
  DFF_X2 \delay1_reg[30]  ( .D(adder_out7[6]), .CK(clock), .Q(delay1[30]) );
  DFF_X2 \delay1_reg[31]  ( .D(adder_out7[7]), .CK(clock), .Q(delay1[31]) );
  DFF_X2 \delay1_reg[32]  ( .D(adder_out7[8]), .CK(clock), .Q(delay1[32]) );
  DFF_X2 \delay1_reg[33]  ( .D(adder_out7[9]), .CK(clock), .Q(delay1[33]) );
  DFF_X2 \delay1_reg[34]  ( .D(adder_out7[10]), .CK(clock), .Q(delay1[34]) );
  DFF_X2 \delay1_reg[35]  ( .D(adder_out7[11]), .CK(clock), .Q(delay1[35]) );
  DFF_X2 \delay1_reg[36]  ( .D(adder_out7[12]), .CK(clock), .Q(delay1[36]) );
  DFF_X2 \delay1_reg[37]  ( .D(adder_out7[13]), .CK(clock), .Q(delay1[37]) );
  DFF_X2 \delay1_reg[38]  ( .D(adder_out7[14]), .CK(clock), .Q(delay1[38]) );
  DFF_X2 \delay1_reg[39]  ( .D(adder_out7[15]), .CK(clock), .Q(delay1[39]) );
  DFF_X2 \delay1_reg[40]  ( .D(adder_out7[16]), .CK(clock), .Q(delay1[40]) );
  DFF_X2 \delay1_reg[41]  ( .D(adder_out7[17]), .CK(clock), .Q(delay1[41]) );
  DFF_X2 \delay1_reg[42]  ( .D(adder_out7[18]), .CK(clock), .Q(delay1[42]) );
  DFF_X2 \delay1_reg[43]  ( .D(adder_out7[19]), .CK(clock), .Q(delay1[43]) );
  DFF_X2 \delay1_reg[44]  ( .D(adder_out7[20]), .CK(clock), .Q(delay1[44]) );
  DFF_X2 \delay1_reg[45]  ( .D(adder_out7[21]), .CK(clock), .Q(delay1[45]) );
  DFF_X2 \delay1_reg[46]  ( .D(adder_out7[22]), .CK(clock), .Q(delay1[46]) );
  DFF_X2 \delay1_reg[47]  ( .D(adder_out7[23]), .CK(clock), .Q(delay1[47]) );
  DFF_X2 \d19_reg[0]  ( .D(d18[0]), .CK(clock), .Q(Mul_In[0]) );
  DFF_X2 \d19_reg[1]  ( .D(d18[1]), .CK(clock), .Q(Mul_In[1]) );
  DFF_X2 \d19_reg[2]  ( .D(d18[2]), .CK(clock), .Q(Mul_In[2]) );
  DFF_X2 \d19_reg[3]  ( .D(d18[3]), .CK(clock), .Q(Mul_In[3]) );
  DFF_X2 \d19_reg[4]  ( .D(d18[4]), .CK(clock), .Q(Mul_In[4]) );
  DFF_X2 \d19_reg[5]  ( .D(d18[5]), .CK(clock), .Q(Mul_In[5]) );
  DFF_X2 \d19_reg[6]  ( .D(d18[6]), .CK(clock), .Q(Mul_In[6]) );
  DFF_X2 \d19_reg[7]  ( .D(d18[7]), .CK(clock), .Q(Mul_In[7]) );
  DFF_X2 \d19_reg[8]  ( .D(d18[8]), .CK(clock), .Q(Mul_In[8]) );
  DFF_X2 \d19_reg[9]  ( .D(d18[9]), .CK(clock), .Q(Mul_In[9]) );
  DFF_X2 \d19_reg[10]  ( .D(d18[10]), .CK(clock), .Q(Mul_In[10]) );
  DFF_X2 \d19_reg[11]  ( .D(d18[11]), .CK(clock), .Q(Mul_In[11]) );
  DFF_X2 \d19_reg[12]  ( .D(d18[12]), .CK(clock), .Q(Mul_In[12]) );
  DFF_X2 \d19_reg[13]  ( .D(d18[13]), .CK(clock), .Q(Mul_In[13]) );
  DFF_X2 \d19_reg[14]  ( .D(d18[14]), .CK(clock), .Q(Mul_In[14]) );
  DFF_X2 \d19_reg[15]  ( .D(d18[15]), .CK(clock), .Q(Mul_In[15]) );
  DFF_X2 \d19_reg[16]  ( .D(d18[16]), .CK(clock), .Q(Mul_In[16]) );
  DFF_X2 \d19_reg[17]  ( .D(d18[17]), .CK(clock), .Q(Mul_In[17]) );
  DFF_X2 \d19_reg[18]  ( .D(d18[18]), .CK(clock), .Q(Mul_In[18]) );
  DFF_X2 \d19_reg[19]  ( .D(d18[19]), .CK(clock), .Q(Mul_In[19]) );
  DFF_X2 \d19_reg[20]  ( .D(d18[20]), .CK(clock), .Q(Mul_In[20]) );
  DFF_X2 \d19_reg[21]  ( .D(d18[21]), .CK(clock), .Q(Mul_In[21]) );
  DFF_X2 \d19_reg[22]  ( .D(d18[22]), .CK(clock), .Q(Mul_In[22]) );
  DFF_X2 \d19_reg[23]  ( .D(d18[23]), .CK(clock), .Q(Mul_In[23]) );
  DFF_X2 \d19_reg[24]  ( .D(d18[24]), .CK(clock), .Q(Mul_In[24]) );
  DFF_X2 \d19_reg[25]  ( .D(d18[25]), .CK(clock), .Q(Mul_In[25]) );
  DFF_X2 \d19_reg[26]  ( .D(d18[26]), .CK(clock), .Q(Mul_In[26]) );
  DFF_X2 \d19_reg[27]  ( .D(d18[27]), .CK(clock), .Q(Mul_In[27]) );
  DFF_X2 \d19_reg[28]  ( .D(d18[28]), .CK(clock), .Q(Mul_In[28]) );
  DFF_X2 \d19_reg[29]  ( .D(d18[29]), .CK(clock), .Q(Mul_In[29]) );
  DFF_X2 \d19_reg[30]  ( .D(d18[30]), .CK(clock), .Q(Mul_In[30]) );
  DFF_X2 \d19_reg[31]  ( .D(d18[31]), .CK(clock), .Q(Mul_In[31]) );
  DFF_X2 \d19_reg[32]  ( .D(d18[32]), .CK(clock), .Q(Mul_In[32]) );
  DFF_X2 \d19_reg[33]  ( .D(d18[33]), .CK(clock), .Q(Mul_In[33]) );
  DFF_X2 \d19_reg[34]  ( .D(d18[34]), .CK(clock), .Q(Mul_In[34]) );
  DFF_X2 \d19_reg[35]  ( .D(d18[35]), .CK(clock), .Q(Mul_In[35]) );
  DFF_X2 \d19_reg[36]  ( .D(d18[36]), .CK(clock), .Q(Mul_In[36]) );
  DFF_X2 \d19_reg[37]  ( .D(d18[37]), .CK(clock), .Q(Mul_In[37]) );
  DFF_X2 \d19_reg[38]  ( .D(d18[38]), .CK(clock), .Q(Mul_In[38]) );
  DFF_X2 \d19_reg[39]  ( .D(d18[39]), .CK(clock), .Q(Mul_In[39]) );
  DFF_X2 \d19_reg[40]  ( .D(d18[40]), .CK(clock), .Q(Mul_In[40]) );
  DFF_X2 \d19_reg[41]  ( .D(d18[41]), .CK(clock), .Q(Mul_In[41]) );
  DFF_X2 \d19_reg[42]  ( .D(d18[42]), .CK(clock), .Q(Mul_In[42]) );
  DFF_X2 \d19_reg[43]  ( .D(d18[43]), .CK(clock), .Q(Mul_In[43]) );
  DFF_X2 \d19_reg[44]  ( .D(d18[44]), .CK(clock), .Q(Mul_In[44]) );
  DFF_X2 \d19_reg[45]  ( .D(d18[45]), .CK(clock), .Q(Mul_In[45]) );
  DFF_X2 \d19_reg[46]  ( .D(d18[46]), .CK(clock), .Q(Mul_In[46]) );
  DFF_X2 \d19_reg[47]  ( .D(d18[47]), .CK(clock), .Q(Mul_In[47]) );
  DFF_X2 \op_reg_reg[0]  ( .D(op_final[0]), .CK(clock), .Q(op_reg[0]) );
  DFF_X2 \op_reg_reg[10]  ( .D(op_final[10]), .CK(clock), .Q(op_reg[10]) );
  DFF_X2 \op_reg_reg[2]  ( .D(op_final[2]), .CK(clock), .Q(op_reg[2]) );
  DFF_X2 \op_reg_reg[6]  ( .D(op_final[6]), .CK(clock), .Q(op_reg[6]) );
  DFF_X2 \op_reg_reg[35]  ( .D(op_final[35]), .CK(clock), .Q(op_reg[35]) );
  DFF_X2 \op_reg_reg[13]  ( .D(op_final[13]), .CK(clock), .Q(op_reg[13]) );
  DFF_X2 \op_reg_reg[21]  ( .D(op_final[21]), .CK(clock), .Q(op_reg[21]) );
  DFF_X2 \op_reg_reg[32]  ( .D(op_final[32]), .CK(clock), .Q(op_reg[32]) );
  DFF_X2 \op_reg_reg[43]  ( .D(op_final[43]), .CK(clock), .Q(op_reg[43]) );
  DFF_X2 \op_reg_reg[16]  ( .D(op_final[16]), .CK(clock), .Q(op_reg[16]) );
  DFF_X2 \op_reg_reg[9]  ( .D(op_final[9]), .CK(clock), .Q(op_reg[9]) );
  DFF_X2 \op_reg_reg[24]  ( .D(op_final[24]), .CK(clock), .Q(op_reg[24]) );
  DFF_X2 \op_reg_reg[38]  ( .D(op_final[38]), .CK(clock), .Q(op_reg[38]) );
  DFF_X2 \op_reg_reg[19]  ( .D(op_final[19]), .CK(clock), .Q(op_reg[19]) );
  DFF_X2 \op_reg_reg[27]  ( .D(op_final[27]), .CK(clock), .Q(op_reg[27]) );
  DFF_X2 \op_reg_reg[40]  ( .D(op_final[40]), .CK(clock), .Q(op_reg[40]) );
  DFF_X2 \op_reg_reg[46]  ( .D(op_final[46]), .CK(clock), .Q(op_reg[46]) );
  DFF_X2 \op_reg_reg[18]  ( .D(op_final[18]), .CK(clock), .Q(op_reg[18]) );
  DFF_X2 \op_reg_reg[8]  ( .D(op_final[8]), .CK(clock), .Q(op_reg[8]) );
  DFF_X2 \op_reg_reg[26]  ( .D(op_final[26]), .CK(clock), .Q(op_reg[26]) );
  DFF_X2 \op_reg_reg[34]  ( .D(op_final[34]), .CK(clock), .Q(op_reg[34]) );
  DFF_X2 \op_reg_reg[29]  ( .D(op_final[29]), .CK(clock), .Q(op_reg[29]) );
  DFF_X2 \op_reg_reg[37]  ( .D(op_final[37]), .CK(clock), .Q(op_reg[37]) );
  DFF_X2 \op_reg_reg[45]  ( .D(op_final[45]), .CK(clock), .Q(op_reg[45]) );
  INV_X4 U52 ( .A(1'b1), .ZN(adder_out4_imag[0]) );
  INV_X4 U54 ( .A(1'b1), .ZN(adder_out4_imag[1]) );
  INV_X4 U56 ( .A(1'b1), .ZN(adder_out4_imag[2]) );
  INV_X4 U58 ( .A(1'b1), .ZN(adder_out4_imag[3]) );
  INV_X4 U60 ( .A(1'b1), .ZN(adder_out4_imag[4]) );
  INV_X4 U62 ( .A(1'b1), .ZN(adder_out4_imag[5]) );
  INV_X4 U64 ( .A(1'b1), .ZN(adder_out4_imag[6]) );
  INV_X4 U66 ( .A(1'b1), .ZN(adder_out4_imag[7]) );
  INV_X4 U68 ( .A(1'b1), .ZN(adder_out4_imag[8]) );
  INV_X4 U70 ( .A(1'b1), .ZN(adder_out4_imag[9]) );
  INV_X4 U72 ( .A(1'b1), .ZN(adder_out4_imag[10]) );
  INV_X4 U74 ( .A(1'b1), .ZN(adder_out4_imag[11]) );
  INV_X4 U76 ( .A(1'b1), .ZN(adder_out4_imag[12]) );
  INV_X4 U78 ( .A(1'b1), .ZN(adder_out4_imag[13]) );
  INV_X4 U80 ( .A(1'b1), .ZN(adder_out4_imag[14]) );
  INV_X4 U82 ( .A(1'b1), .ZN(adder_out4_imag[15]) );
  INV_X4 U84 ( .A(1'b1), .ZN(adder_out4_imag[16]) );
  INV_X4 U86 ( .A(1'b1), .ZN(adder_out4_imag[17]) );
  INV_X4 U88 ( .A(1'b1), .ZN(adder_out4_imag[18]) );
  INV_X4 U90 ( .A(1'b1), .ZN(adder_out4_imag[19]) );
  INV_X4 U92 ( .A(1'b1), .ZN(adder_out4_imag[20]) );
  INV_X4 U94 ( .A(1'b1), .ZN(adder_out4_imag[21]) );
  INV_X4 U96 ( .A(1'b1), .ZN(adder_out4_imag[22]) );
  INV_X4 U98 ( .A(1'b1), .ZN(adder_out4_imag[23]) );
  INV_X4 U100 ( .A(1'b1), .ZN(adder_out3_imag[0]) );
  INV_X4 U102 ( .A(1'b1), .ZN(adder_out3_imag[1]) );
  INV_X4 U104 ( .A(1'b1), .ZN(adder_out3_imag[2]) );
  INV_X4 U106 ( .A(1'b1), .ZN(adder_out3_imag[3]) );
  INV_X4 U108 ( .A(1'b1), .ZN(adder_out3_imag[4]) );
  INV_X4 U110 ( .A(1'b1), .ZN(adder_out3_imag[5]) );
  INV_X4 U112 ( .A(1'b1), .ZN(adder_out3_imag[6]) );
  INV_X4 U114 ( .A(1'b1), .ZN(adder_out3_imag[7]) );
  INV_X4 U116 ( .A(1'b1), .ZN(adder_out3_imag[8]) );
  INV_X4 U118 ( .A(1'b1), .ZN(adder_out3_imag[9]) );
  INV_X4 U120 ( .A(1'b1), .ZN(adder_out3_imag[10]) );
  INV_X4 U122 ( .A(1'b1), .ZN(adder_out3_imag[11]) );
  INV_X4 U124 ( .A(1'b1), .ZN(adder_out3_imag[12]) );
  INV_X4 U126 ( .A(1'b1), .ZN(adder_out3_imag[13]) );
  INV_X4 U128 ( .A(1'b1), .ZN(adder_out3_imag[14]) );
  INV_X4 U130 ( .A(1'b1), .ZN(adder_out3_imag[15]) );
  INV_X4 U132 ( .A(1'b1), .ZN(adder_out3_imag[16]) );
  INV_X4 U134 ( .A(1'b1), .ZN(adder_out3_imag[17]) );
  INV_X4 U136 ( .A(1'b1), .ZN(adder_out3_imag[18]) );
  INV_X4 U138 ( .A(1'b1), .ZN(adder_out3_imag[19]) );
  INV_X4 U140 ( .A(1'b1), .ZN(adder_out3_imag[20]) );
  INV_X4 U142 ( .A(1'b1), .ZN(adder_out3_imag[21]) );
  INV_X4 U144 ( .A(1'b1), .ZN(adder_out3_imag[22]) );
  INV_X4 U146 ( .A(1'b1), .ZN(adder_out3_imag[23]) );
  INV_X4 U148 ( .A(1'b1), .ZN(adder_out4[0]) );
  INV_X4 U150 ( .A(1'b1), .ZN(adder_out4[1]) );
  INV_X4 U152 ( .A(1'b1), .ZN(adder_out4[2]) );
  INV_X4 U154 ( .A(1'b1), .ZN(adder_out4[3]) );
  INV_X4 U156 ( .A(1'b1), .ZN(adder_out4[4]) );
  INV_X4 U158 ( .A(1'b1), .ZN(adder_out4[5]) );
  INV_X4 U160 ( .A(1'b1), .ZN(adder_out4[6]) );
  INV_X4 U162 ( .A(1'b1), .ZN(adder_out4[7]) );
  INV_X4 U164 ( .A(1'b1), .ZN(adder_out4[8]) );
  INV_X4 U166 ( .A(1'b1), .ZN(adder_out4[9]) );
  INV_X4 U168 ( .A(1'b1), .ZN(adder_out4[10]) );
  INV_X4 U170 ( .A(1'b1), .ZN(adder_out4[11]) );
  INV_X4 U172 ( .A(1'b1), .ZN(adder_out4[12]) );
  INV_X4 U174 ( .A(1'b1), .ZN(adder_out4[13]) );
  INV_X4 U176 ( .A(1'b1), .ZN(adder_out4[14]) );
  INV_X4 U178 ( .A(1'b1), .ZN(adder_out4[15]) );
  INV_X4 U180 ( .A(1'b1), .ZN(adder_out4[16]) );
  INV_X4 U182 ( .A(1'b1), .ZN(adder_out4[17]) );
  INV_X4 U184 ( .A(1'b1), .ZN(adder_out4[18]) );
  INV_X4 U186 ( .A(1'b1), .ZN(adder_out4[19]) );
  INV_X4 U188 ( .A(1'b1), .ZN(adder_out4[20]) );
  INV_X4 U190 ( .A(1'b1), .ZN(adder_out4[21]) );
  INV_X4 U192 ( .A(1'b1), .ZN(adder_out4[22]) );
  INV_X4 U194 ( .A(1'b1), .ZN(adder_out4[23]) );
  INV_X4 U196 ( .A(1'b1), .ZN(adder_out3[0]) );
  INV_X4 U198 ( .A(1'b1), .ZN(adder_out3[1]) );
  INV_X4 U200 ( .A(1'b1), .ZN(adder_out3[2]) );
  INV_X4 U202 ( .A(1'b1), .ZN(adder_out3[3]) );
  INV_X4 U204 ( .A(1'b1), .ZN(adder_out3[4]) );
  INV_X4 U206 ( .A(1'b1), .ZN(adder_out3[5]) );
  INV_X4 U208 ( .A(1'b1), .ZN(adder_out3[6]) );
  INV_X4 U210 ( .A(1'b1), .ZN(adder_out3[7]) );
  INV_X4 U212 ( .A(1'b1), .ZN(adder_out3[8]) );
  INV_X4 U214 ( .A(1'b1), .ZN(adder_out3[9]) );
  INV_X4 U216 ( .A(1'b1), .ZN(adder_out3[10]) );
  INV_X4 U218 ( .A(1'b1), .ZN(adder_out3[11]) );
  INV_X4 U220 ( .A(1'b1), .ZN(adder_out3[12]) );
  INV_X4 U222 ( .A(1'b1), .ZN(adder_out3[13]) );
  INV_X4 U224 ( .A(1'b1), .ZN(adder_out3[14]) );
  INV_X4 U226 ( .A(1'b1), .ZN(adder_out3[15]) );
  INV_X4 U228 ( .A(1'b1), .ZN(adder_out3[16]) );
  INV_X4 U230 ( .A(1'b1), .ZN(adder_out3[17]) );
  INV_X4 U232 ( .A(1'b1), .ZN(adder_out3[18]) );
  INV_X4 U234 ( .A(1'b1), .ZN(adder_out3[19]) );
  INV_X4 U236 ( .A(1'b1), .ZN(adder_out3[20]) );
  INV_X4 U238 ( .A(1'b1), .ZN(adder_out3[21]) );
  INV_X4 U240 ( .A(1'b1), .ZN(adder_out3[22]) );
  INV_X4 U242 ( .A(1'b1), .ZN(adder_out3[23]) );
  INV_X4 U244 ( .A(1'b1), .ZN(adder_out2_imag[0]) );
  INV_X4 U246 ( .A(1'b1), .ZN(adder_out2_imag[1]) );
  INV_X4 U248 ( .A(1'b1), .ZN(adder_out2_imag[2]) );
  INV_X4 U250 ( .A(1'b1), .ZN(adder_out2_imag[3]) );
  INV_X4 U252 ( .A(1'b1), .ZN(adder_out2_imag[4]) );
  INV_X4 U254 ( .A(1'b1), .ZN(adder_out2_imag[5]) );
  INV_X4 U256 ( .A(1'b1), .ZN(adder_out2_imag[6]) );
  INV_X4 U258 ( .A(1'b1), .ZN(adder_out2_imag[7]) );
  INV_X4 U260 ( .A(1'b1), .ZN(adder_out2_imag[8]) );
  INV_X4 U262 ( .A(1'b1), .ZN(adder_out2_imag[9]) );
  INV_X4 U264 ( .A(1'b1), .ZN(adder_out2_imag[10]) );
  INV_X4 U266 ( .A(1'b1), .ZN(adder_out2_imag[11]) );
  INV_X4 U268 ( .A(1'b1), .ZN(adder_out2_imag[12]) );
  INV_X4 U270 ( .A(1'b1), .ZN(adder_out2_imag[13]) );
  INV_X4 U272 ( .A(1'b1), .ZN(adder_out2_imag[14]) );
  INV_X4 U274 ( .A(1'b1), .ZN(adder_out2_imag[15]) );
  INV_X4 U276 ( .A(1'b1), .ZN(adder_out2_imag[16]) );
  INV_X4 U278 ( .A(1'b1), .ZN(adder_out2_imag[17]) );
  INV_X4 U280 ( .A(1'b1), .ZN(adder_out2_imag[18]) );
  INV_X4 U282 ( .A(1'b1), .ZN(adder_out2_imag[19]) );
  INV_X4 U284 ( .A(1'b1), .ZN(adder_out2_imag[20]) );
  INV_X4 U286 ( .A(1'b1), .ZN(adder_out2_imag[21]) );
  INV_X4 U288 ( .A(1'b1), .ZN(adder_out2_imag[22]) );
  INV_X4 U290 ( .A(1'b1), .ZN(adder_out2_imag[23]) );
  INV_X4 U292 ( .A(1'b1), .ZN(adder_out1_imag[0]) );
  INV_X4 U294 ( .A(1'b1), .ZN(adder_out1_imag[1]) );
  INV_X4 U296 ( .A(1'b1), .ZN(adder_out1_imag[2]) );
  INV_X4 U298 ( .A(1'b1), .ZN(adder_out1_imag[3]) );
  INV_X4 U300 ( .A(1'b1), .ZN(adder_out1_imag[4]) );
  INV_X4 U302 ( .A(1'b1), .ZN(adder_out1_imag[5]) );
  INV_X4 U304 ( .A(1'b1), .ZN(adder_out1_imag[6]) );
  INV_X4 U306 ( .A(1'b1), .ZN(adder_out1_imag[7]) );
  INV_X4 U308 ( .A(1'b1), .ZN(adder_out1_imag[8]) );
  INV_X4 U310 ( .A(1'b1), .ZN(adder_out1_imag[9]) );
  INV_X4 U312 ( .A(1'b1), .ZN(adder_out1_imag[10]) );
  INV_X4 U314 ( .A(1'b1), .ZN(adder_out1_imag[11]) );
  INV_X4 U316 ( .A(1'b1), .ZN(adder_out1_imag[12]) );
  INV_X4 U318 ( .A(1'b1), .ZN(adder_out1_imag[13]) );
  INV_X4 U320 ( .A(1'b1), .ZN(adder_out1_imag[14]) );
  INV_X4 U322 ( .A(1'b1), .ZN(adder_out1_imag[15]) );
  INV_X4 U324 ( .A(1'b1), .ZN(adder_out1_imag[16]) );
  INV_X4 U326 ( .A(1'b1), .ZN(adder_out1_imag[17]) );
  INV_X4 U328 ( .A(1'b1), .ZN(adder_out1_imag[18]) );
  INV_X4 U330 ( .A(1'b1), .ZN(adder_out1_imag[19]) );
  INV_X4 U332 ( .A(1'b1), .ZN(adder_out1_imag[20]) );
  INV_X4 U334 ( .A(1'b1), .ZN(adder_out1_imag[21]) );
  INV_X4 U336 ( .A(1'b1), .ZN(adder_out1_imag[22]) );
  INV_X4 U338 ( .A(1'b1), .ZN(adder_out1_imag[23]) );
  INV_X4 U340 ( .A(1'b1), .ZN(adder_out2[0]) );
  INV_X4 U342 ( .A(1'b1), .ZN(adder_out2[1]) );
  INV_X4 U344 ( .A(1'b1), .ZN(adder_out2[2]) );
  INV_X4 U346 ( .A(1'b1), .ZN(adder_out2[3]) );
  INV_X4 U348 ( .A(1'b1), .ZN(adder_out2[4]) );
  INV_X4 U350 ( .A(1'b1), .ZN(adder_out2[5]) );
  INV_X4 U352 ( .A(1'b1), .ZN(adder_out2[6]) );
  INV_X4 U354 ( .A(1'b1), .ZN(adder_out2[7]) );
  INV_X4 U356 ( .A(1'b1), .ZN(adder_out2[8]) );
  INV_X4 U358 ( .A(1'b1), .ZN(adder_out2[9]) );
  INV_X4 U360 ( .A(1'b1), .ZN(adder_out2[10]) );
  INV_X4 U362 ( .A(1'b1), .ZN(adder_out2[11]) );
  INV_X4 U364 ( .A(1'b1), .ZN(adder_out2[12]) );
  INV_X4 U366 ( .A(1'b1), .ZN(adder_out2[13]) );
  INV_X4 U368 ( .A(1'b1), .ZN(adder_out2[14]) );
  INV_X4 U370 ( .A(1'b1), .ZN(adder_out2[15]) );
  INV_X4 U372 ( .A(1'b1), .ZN(adder_out2[16]) );
  INV_X4 U374 ( .A(1'b1), .ZN(adder_out2[17]) );
  INV_X4 U376 ( .A(1'b1), .ZN(adder_out2[18]) );
  INV_X4 U378 ( .A(1'b1), .ZN(adder_out2[19]) );
  INV_X4 U380 ( .A(1'b1), .ZN(adder_out2[20]) );
  INV_X4 U382 ( .A(1'b1), .ZN(adder_out2[21]) );
  INV_X4 U384 ( .A(1'b1), .ZN(adder_out2[22]) );
  INV_X4 U386 ( .A(1'b1), .ZN(adder_out2[23]) );
  INV_X4 U388 ( .A(1'b1), .ZN(adder_out1[0]) );
  INV_X4 U390 ( .A(1'b1), .ZN(adder_out1[1]) );
  INV_X4 U392 ( .A(1'b1), .ZN(adder_out1[2]) );
  INV_X4 U394 ( .A(1'b1), .ZN(adder_out1[3]) );
  INV_X4 U396 ( .A(1'b1), .ZN(adder_out1[4]) );
  INV_X4 U398 ( .A(1'b1), .ZN(adder_out1[5]) );
  INV_X4 U400 ( .A(1'b1), .ZN(adder_out1[6]) );
  INV_X4 U402 ( .A(1'b1), .ZN(adder_out1[7]) );
  INV_X4 U404 ( .A(1'b1), .ZN(adder_out1[8]) );
  INV_X4 U406 ( .A(1'b1), .ZN(adder_out1[9]) );
  INV_X4 U408 ( .A(1'b1), .ZN(adder_out1[10]) );
  INV_X4 U410 ( .A(1'b1), .ZN(adder_out1[11]) );
  INV_X4 U412 ( .A(1'b1), .ZN(adder_out1[12]) );
  INV_X4 U414 ( .A(1'b1), .ZN(adder_out1[13]) );
  INV_X4 U416 ( .A(1'b1), .ZN(adder_out1[14]) );
  INV_X4 U418 ( .A(1'b1), .ZN(adder_out1[15]) );
  INV_X4 U420 ( .A(1'b1), .ZN(adder_out1[16]) );
  INV_X4 U422 ( .A(1'b1), .ZN(adder_out1[17]) );
  INV_X4 U424 ( .A(1'b1), .ZN(adder_out1[18]) );
  INV_X4 U426 ( .A(1'b1), .ZN(adder_out1[19]) );
  INV_X4 U428 ( .A(1'b1), .ZN(adder_out1[20]) );
  INV_X4 U430 ( .A(1'b1), .ZN(adder_out1[21]) );
  INV_X4 U432 ( .A(1'b1), .ZN(adder_out1[22]) );
  INV_X4 U434 ( .A(1'b1), .ZN(adder_out1[23]) );
  INV_X4 U436 ( .A(adder_output[24]), .ZN(n903) );
  INV_X4 U437 ( .A(n903), .ZN(n902) );
  INV_X4 U438 ( .A(n688), .ZN(n689) );
  INV_X4 U439 ( .A(ReadBus1[118]), .ZN(n688) );
  INV_X4 U440 ( .A(n696), .ZN(n697) );
  INV_X4 U441 ( .A(ReadBus1[122]), .ZN(n696) );
  INV_X4 U442 ( .A(n704), .ZN(n705) );
  INV_X4 U443 ( .A(ReadBus1[126]), .ZN(n704) );
  INV_X4 U444 ( .A(n706), .ZN(n707) );
  INV_X4 U445 ( .A(ReadBus1[127]), .ZN(n706) );
  INV_X4 U446 ( .A(n580), .ZN(n581) );
  INV_X4 U447 ( .A(ReadBus1[49]), .ZN(n580) );
  INV_X4 U448 ( .A(n582), .ZN(n583) );
  INV_X4 U449 ( .A(ReadBus1[50]), .ZN(n582) );
  INV_X4 U450 ( .A(n680), .ZN(n681) );
  INV_X4 U451 ( .A(ReadBus1[114]), .ZN(n680) );
  INV_X4 U452 ( .A(n584), .ZN(n585) );
  INV_X4 U453 ( .A(ReadBus1[51]), .ZN(n584) );
  INV_X4 U454 ( .A(n682), .ZN(n683) );
  INV_X4 U455 ( .A(ReadBus1[115]), .ZN(n682) );
  INV_X4 U456 ( .A(n588), .ZN(n589) );
  INV_X4 U457 ( .A(ReadBus1[53]), .ZN(n588) );
  INV_X4 U458 ( .A(n590), .ZN(n591) );
  INV_X4 U459 ( .A(ReadBus1[54]), .ZN(n590) );
  INV_X4 U460 ( .A(n592), .ZN(n593) );
  INV_X4 U461 ( .A(ReadBus1[55]), .ZN(n592) );
  INV_X4 U462 ( .A(n690), .ZN(n691) );
  INV_X4 U463 ( .A(ReadBus1[119]), .ZN(n690) );
  INV_X4 U464 ( .A(n598), .ZN(n599) );
  INV_X4 U465 ( .A(ReadBus1[58]), .ZN(n598) );
  INV_X4 U466 ( .A(n596), .ZN(n597) );
  INV_X4 U467 ( .A(ReadBus1[57]), .ZN(n596) );
  INV_X4 U468 ( .A(n600), .ZN(n601) );
  INV_X4 U469 ( .A(ReadBus1[59]), .ZN(n600) );
  INV_X4 U470 ( .A(n604), .ZN(n605) );
  INV_X4 U471 ( .A(ReadBus1[61]), .ZN(n604) );
  INV_X4 U472 ( .A(n606), .ZN(n607) );
  INV_X4 U473 ( .A(ReadBus1[62]), .ZN(n606) );
  INV_X4 U474 ( .A(n608), .ZN(n609) );
  INV_X4 U475 ( .A(ReadBus1[63]), .ZN(n608) );
  INV_X4 U476 ( .A(n698), .ZN(n699) );
  INV_X4 U477 ( .A(ReadBus1[123]), .ZN(n698) );
  INV_X4 U478 ( .A(n772), .ZN(n773) );
  INV_X4 U479 ( .A(Y[0]), .ZN(n772) );
  INV_X4 U480 ( .A(n578), .ZN(n579) );
  INV_X4 U481 ( .A(ReadBus1[48]), .ZN(n578) );
  INV_X4 U482 ( .A(n676), .ZN(n677) );
  INV_X4 U483 ( .A(ReadBus1[112]), .ZN(n676) );
  INV_X4 U484 ( .A(n708), .ZN(n709) );
  INV_X4 U485 ( .A(ReadBus1[176]), .ZN(n708) );
  INV_X4 U486 ( .A(n678), .ZN(n679) );
  INV_X4 U487 ( .A(ReadBus1[113]), .ZN(n678) );
  INV_X4 U488 ( .A(n710), .ZN(n711) );
  INV_X4 U489 ( .A(ReadBus1[177]), .ZN(n710) );
  INV_X4 U490 ( .A(n712), .ZN(n713) );
  INV_X4 U491 ( .A(ReadBus1[178]), .ZN(n712) );
  INV_X4 U492 ( .A(n714), .ZN(n715) );
  INV_X4 U493 ( .A(ReadBus1[179]), .ZN(n714) );
  INV_X4 U494 ( .A(n586), .ZN(n587) );
  INV_X4 U495 ( .A(ReadBus1[52]), .ZN(n586) );
  INV_X4 U496 ( .A(n684), .ZN(n685) );
  INV_X4 U497 ( .A(ReadBus1[116]), .ZN(n684) );
  INV_X4 U498 ( .A(n716), .ZN(n717) );
  INV_X4 U499 ( .A(ReadBus1[180]), .ZN(n716) );
  INV_X4 U500 ( .A(n686), .ZN(n687) );
  INV_X4 U501 ( .A(ReadBus1[117]), .ZN(n686) );
  INV_X4 U502 ( .A(n718), .ZN(n719) );
  INV_X4 U503 ( .A(ReadBus1[181]), .ZN(n718) );
  INV_X4 U504 ( .A(n720), .ZN(n721) );
  INV_X4 U505 ( .A(ReadBus1[182]), .ZN(n720) );
  INV_X4 U506 ( .A(n722), .ZN(n723) );
  INV_X4 U507 ( .A(ReadBus1[183]), .ZN(n722) );
  INV_X4 U508 ( .A(n594), .ZN(n595) );
  INV_X4 U509 ( .A(ReadBus1[56]), .ZN(n594) );
  INV_X4 U510 ( .A(n724), .ZN(n725) );
  INV_X4 U511 ( .A(ReadBus1[184]), .ZN(n724) );
  INV_X4 U512 ( .A(n692), .ZN(n693) );
  INV_X4 U513 ( .A(ReadBus1[120]), .ZN(n692) );
  INV_X4 U514 ( .A(n726), .ZN(n727) );
  INV_X4 U515 ( .A(ReadBus1[185]), .ZN(n726) );
  INV_X4 U516 ( .A(n694), .ZN(n695) );
  INV_X4 U517 ( .A(ReadBus1[121]), .ZN(n694) );
  INV_X4 U518 ( .A(n728), .ZN(n729) );
  INV_X4 U519 ( .A(ReadBus1[186]), .ZN(n728) );
  INV_X4 U520 ( .A(n602), .ZN(n603) );
  INV_X4 U521 ( .A(ReadBus1[60]), .ZN(n602) );
  INV_X4 U522 ( .A(n700), .ZN(n701) );
  INV_X4 U523 ( .A(ReadBus1[124]), .ZN(n700) );
  INV_X4 U524 ( .A(n702), .ZN(n703) );
  INV_X4 U525 ( .A(ReadBus1[125]), .ZN(n702) );
  INV_X4 U526 ( .A(n730), .ZN(n731) );
  INV_X4 U527 ( .A(ReadBus1[187]), .ZN(n730) );
  INV_X4 U528 ( .A(n732), .ZN(n733) );
  INV_X4 U529 ( .A(ReadBus1[188]), .ZN(n732) );
  INV_X4 U530 ( .A(n734), .ZN(n735) );
  INV_X4 U531 ( .A(ReadBus1[189]), .ZN(n734) );
  INV_X4 U532 ( .A(n736), .ZN(n737) );
  INV_X4 U533 ( .A(ReadBus1[190]), .ZN(n736) );
  INV_X4 U534 ( .A(n738), .ZN(n739) );
  INV_X4 U535 ( .A(ReadBus1[191]), .ZN(n738) );
  INV_X4 U536 ( .A(n778), .ZN(n779) );
  INV_X4 U537 ( .A(Y[3]), .ZN(n778) );
  INV_X4 U538 ( .A(n774), .ZN(n775) );
  INV_X4 U539 ( .A(Y[1]), .ZN(n774) );
  INV_X4 U540 ( .A(n776), .ZN(n777) );
  INV_X4 U541 ( .A(Y[2]), .ZN(n776) );
  INV_X4 U542 ( .A(n782), .ZN(n783) );
  INV_X4 U543 ( .A(Y[5]), .ZN(n782) );
  INV_X4 U544 ( .A(n780), .ZN(n781) );
  INV_X4 U545 ( .A(Y[4]), .ZN(n780) );
  INV_X4 U546 ( .A(n784), .ZN(n785) );
  INV_X4 U547 ( .A(Y[6]), .ZN(n784) );
  INV_X4 U548 ( .A(n786), .ZN(n787) );
  INV_X4 U549 ( .A(Y[7]), .ZN(n786) );
  INV_X4 U550 ( .A(n788), .ZN(n789) );
  INV_X4 U551 ( .A(X[0]), .ZN(n788) );
  INV_X4 U552 ( .A(n610), .ZN(n611) );
  INV_X4 U553 ( .A(ReadBus1[64]), .ZN(n610) );
  INV_X4 U554 ( .A(n612), .ZN(n613) );
  INV_X4 U555 ( .A(ReadBus1[65]), .ZN(n612) );
  INV_X4 U556 ( .A(n614), .ZN(n615) );
  INV_X4 U557 ( .A(ReadBus1[66]), .ZN(n614) );
  INV_X4 U558 ( .A(n616), .ZN(n617) );
  INV_X4 U559 ( .A(ReadBus1[67]), .ZN(n616) );
  INV_X4 U560 ( .A(n618), .ZN(n619) );
  INV_X4 U561 ( .A(ReadBus1[68]), .ZN(n618) );
  INV_X4 U562 ( .A(n620), .ZN(n621) );
  INV_X4 U563 ( .A(ReadBus1[69]), .ZN(n620) );
  INV_X4 U564 ( .A(n622), .ZN(n623) );
  INV_X4 U565 ( .A(ReadBus1[70]), .ZN(n622) );
  INV_X4 U566 ( .A(n624), .ZN(n625) );
  INV_X4 U567 ( .A(ReadBus1[71]), .ZN(n624) );
  INV_X4 U568 ( .A(n626), .ZN(n627) );
  INV_X4 U569 ( .A(ReadBus1[72]), .ZN(n626) );
  INV_X4 U570 ( .A(n628), .ZN(n629) );
  INV_X4 U571 ( .A(ReadBus1[73]), .ZN(n628) );
  INV_X4 U572 ( .A(n630), .ZN(n631) );
  INV_X4 U573 ( .A(ReadBus1[74]), .ZN(n630) );
  INV_X4 U574 ( .A(n632), .ZN(n633) );
  INV_X4 U575 ( .A(ReadBus1[80]), .ZN(n632) );
  INV_X4 U576 ( .A(n634), .ZN(n635) );
  INV_X4 U577 ( .A(ReadBus1[81]), .ZN(n634) );
  INV_X4 U578 ( .A(n636), .ZN(n637) );
  INV_X4 U579 ( .A(ReadBus1[82]), .ZN(n636) );
  INV_X4 U580 ( .A(n638), .ZN(n639) );
  INV_X4 U581 ( .A(ReadBus1[83]), .ZN(n638) );
  INV_X4 U582 ( .A(n640), .ZN(n641) );
  INV_X4 U583 ( .A(ReadBus1[84]), .ZN(n640) );
  INV_X4 U584 ( .A(n642), .ZN(n643) );
  INV_X4 U585 ( .A(ReadBus1[85]), .ZN(n642) );
  INV_X4 U586 ( .A(n644), .ZN(n645) );
  INV_X4 U587 ( .A(ReadBus1[86]), .ZN(n644) );
  INV_X4 U588 ( .A(n646), .ZN(n647) );
  INV_X4 U589 ( .A(ReadBus1[87]), .ZN(n646) );
  INV_X4 U590 ( .A(n648), .ZN(n649) );
  INV_X4 U591 ( .A(ReadBus1[88]), .ZN(n648) );
  INV_X4 U592 ( .A(n650), .ZN(n651) );
  INV_X4 U593 ( .A(ReadBus1[89]), .ZN(n650) );
  INV_X4 U594 ( .A(n652), .ZN(n653) );
  INV_X4 U595 ( .A(ReadBus1[90]), .ZN(n652) );
  INV_X4 U596 ( .A(n654), .ZN(n655) );
  INV_X4 U597 ( .A(ReadBus1[96]), .ZN(n654) );
  INV_X4 U598 ( .A(n656), .ZN(n657) );
  INV_X4 U599 ( .A(ReadBus1[97]), .ZN(n656) );
  INV_X4 U600 ( .A(n658), .ZN(n659) );
  INV_X4 U601 ( .A(ReadBus1[98]), .ZN(n658) );
  INV_X4 U602 ( .A(n660), .ZN(n661) );
  INV_X4 U603 ( .A(ReadBus1[99]), .ZN(n660) );
  INV_X4 U604 ( .A(n662), .ZN(n663) );
  INV_X4 U605 ( .A(ReadBus1[100]), .ZN(n662) );
  INV_X4 U606 ( .A(n664), .ZN(n665) );
  INV_X4 U607 ( .A(ReadBus1[101]), .ZN(n664) );
  INV_X4 U608 ( .A(n666), .ZN(n667) );
  INV_X4 U609 ( .A(ReadBus1[102]), .ZN(n666) );
  INV_X4 U610 ( .A(n668), .ZN(n669) );
  INV_X4 U611 ( .A(ReadBus1[103]), .ZN(n668) );
  INV_X4 U612 ( .A(n670), .ZN(n671) );
  INV_X4 U613 ( .A(ReadBus1[104]), .ZN(n670) );
  INV_X4 U614 ( .A(n672), .ZN(n673) );
  INV_X4 U615 ( .A(ReadBus1[105]), .ZN(n672) );
  INV_X4 U616 ( .A(n674), .ZN(n675) );
  INV_X4 U617 ( .A(ReadBus1[106]), .ZN(n674) );
  INV_X4 U618 ( .A(n740), .ZN(n741) );
  INV_X4 U619 ( .A(ReadBus1[240]), .ZN(n740) );
  INV_X4 U620 ( .A(n742), .ZN(n743) );
  INV_X4 U621 ( .A(ReadBus1[241]), .ZN(n742) );
  INV_X4 U622 ( .A(n744), .ZN(n745) );
  INV_X4 U623 ( .A(ReadBus1[242]), .ZN(n744) );
  INV_X4 U624 ( .A(n746), .ZN(n747) );
  INV_X4 U625 ( .A(ReadBus1[243]), .ZN(n746) );
  INV_X4 U626 ( .A(n748), .ZN(n749) );
  INV_X4 U627 ( .A(ReadBus1[244]), .ZN(n748) );
  INV_X4 U628 ( .A(n750), .ZN(n751) );
  INV_X4 U629 ( .A(ReadBus1[245]), .ZN(n750) );
  INV_X4 U630 ( .A(n752), .ZN(n753) );
  INV_X4 U631 ( .A(ReadBus1[246]), .ZN(n752) );
  INV_X4 U632 ( .A(n754), .ZN(n755) );
  INV_X4 U633 ( .A(ReadBus1[247]), .ZN(n754) );
  INV_X4 U634 ( .A(n756), .ZN(n757) );
  INV_X4 U635 ( .A(ReadBus1[248]), .ZN(n756) );
  INV_X4 U636 ( .A(n758), .ZN(n759) );
  INV_X4 U637 ( .A(ReadBus1[249]), .ZN(n758) );
  INV_X4 U638 ( .A(n760), .ZN(n761) );
  INV_X4 U639 ( .A(ReadBus1[250]), .ZN(n760) );
  INV_X4 U640 ( .A(n762), .ZN(n763) );
  INV_X4 U641 ( .A(ReadBus1[251]), .ZN(n762) );
  INV_X4 U642 ( .A(n764), .ZN(n765) );
  INV_X4 U643 ( .A(ReadBus1[252]), .ZN(n764) );
  INV_X4 U644 ( .A(n766), .ZN(n767) );
  INV_X4 U645 ( .A(ReadBus1[253]), .ZN(n766) );
  INV_X4 U646 ( .A(n768), .ZN(n769) );
  INV_X4 U647 ( .A(ReadBus1[254]), .ZN(n768) );
  INV_X4 U648 ( .A(n770), .ZN(n771) );
  INV_X4 U649 ( .A(ReadBus1[255]), .ZN(n770) );
  INV_X4 U650 ( .A(n794), .ZN(n795) );
  INV_X4 U651 ( .A(X[3]), .ZN(n794) );
  INV_X4 U652 ( .A(n790), .ZN(n791) );
  INV_X4 U653 ( .A(X[1]), .ZN(n790) );
  INV_X4 U654 ( .A(n792), .ZN(n793) );
  INV_X4 U655 ( .A(X[2]), .ZN(n792) );
  INV_X4 U656 ( .A(n798), .ZN(n799) );
  INV_X4 U657 ( .A(X[5]), .ZN(n798) );
  INV_X4 U658 ( .A(n796), .ZN(n797) );
  INV_X4 U659 ( .A(X[4]), .ZN(n796) );
  INV_X4 U660 ( .A(n800), .ZN(n801) );
  INV_X4 U661 ( .A(X[6]), .ZN(n800) );
  INV_X4 U662 ( .A(n802), .ZN(n803) );
  INV_X4 U663 ( .A(X[7]), .ZN(n802) );
  INV_X4 U664 ( .A(n816), .ZN(n817) );
  INV_X4 U665 ( .A(multinput[6]), .ZN(n816) );
  INV_X4 U666 ( .A(n864), .ZN(n865) );
  INV_X4 U667 ( .A(multinput[30]), .ZN(n864) );
  INV_X4 U668 ( .A(n866), .ZN(n867) );
  INV_X4 U669 ( .A(multinput[31]), .ZN(n866) );
  INV_X4 U670 ( .A(n868), .ZN(n869) );
  INV_X4 U671 ( .A(multinput[32]), .ZN(n868) );
  INV_X4 U672 ( .A(n822), .ZN(n823) );
  INV_X4 U673 ( .A(multinput[9]), .ZN(n822) );
  INV_X4 U674 ( .A(n812), .ZN(n813) );
  INV_X4 U675 ( .A(multinput[4]), .ZN(n812) );
  INV_X4 U676 ( .A(n824), .ZN(n825) );
  INV_X4 U677 ( .A(multinput[10]), .ZN(n824) );
  INV_X4 U678 ( .A(n830), .ZN(n831) );
  INV_X4 U679 ( .A(multinput[13]), .ZN(n830) );
  INV_X4 U680 ( .A(n836), .ZN(n837) );
  INV_X4 U681 ( .A(multinput[16]), .ZN(n836) );
  INV_X4 U682 ( .A(n842), .ZN(n843) );
  INV_X4 U683 ( .A(multinput[19]), .ZN(n842) );
  INV_X4 U684 ( .A(n846), .ZN(n847) );
  INV_X4 U685 ( .A(multinput[21]), .ZN(n846) );
  INV_X4 U686 ( .A(n872), .ZN(n873) );
  INV_X4 U687 ( .A(multinput[34]), .ZN(n872) );
  INV_X4 U688 ( .A(n878), .ZN(n879) );
  INV_X4 U689 ( .A(multinput[37]), .ZN(n878) );
  INV_X4 U690 ( .A(n884), .ZN(n885) );
  INV_X4 U691 ( .A(multinput[40]), .ZN(n884) );
  INV_X4 U692 ( .A(n890), .ZN(n891) );
  INV_X4 U693 ( .A(multinput[43]), .ZN(n890) );
  INV_X4 U694 ( .A(n806), .ZN(n807) );
  INV_X4 U695 ( .A(multinput[1]), .ZN(n806) );
  INV_X4 U696 ( .A(n808), .ZN(n809) );
  INV_X4 U697 ( .A(multinput[2]), .ZN(n808) );
  INV_X4 U698 ( .A(n814), .ZN(n815) );
  INV_X4 U699 ( .A(multinput[5]), .ZN(n814) );
  INV_X4 U700 ( .A(n826), .ZN(n827) );
  INV_X4 U701 ( .A(multinput[11]), .ZN(n826) );
  INV_X4 U702 ( .A(n832), .ZN(n833) );
  INV_X4 U703 ( .A(multinput[14]), .ZN(n832) );
  INV_X4 U704 ( .A(n838), .ZN(n839) );
  INV_X4 U705 ( .A(multinput[17]), .ZN(n838) );
  INV_X4 U706 ( .A(n848), .ZN(n849) );
  INV_X4 U707 ( .A(multinput[22]), .ZN(n848) );
  INV_X4 U708 ( .A(n900), .ZN(n901) );
  INV_X4 U709 ( .A(reset), .ZN(n900) );
  INV_X4 U710 ( .A(n804), .ZN(n805) );
  INV_X4 U711 ( .A(multinput[0]), .ZN(n804) );
  INV_X4 U712 ( .A(n810), .ZN(n811) );
  INV_X4 U713 ( .A(multinput[3]), .ZN(n810) );
  INV_X4 U714 ( .A(n818), .ZN(n819) );
  INV_X4 U715 ( .A(multinput[7]), .ZN(n818) );
  INV_X4 U716 ( .A(n820), .ZN(n821) );
  INV_X4 U717 ( .A(multinput[8]), .ZN(n820) );
  INV_X4 U718 ( .A(n828), .ZN(n829) );
  INV_X4 U719 ( .A(multinput[12]), .ZN(n828) );
  INV_X4 U720 ( .A(n834), .ZN(n835) );
  INV_X4 U721 ( .A(multinput[15]), .ZN(n834) );
  INV_X4 U722 ( .A(n840), .ZN(n841) );
  INV_X4 U723 ( .A(multinput[18]), .ZN(n840) );
  INV_X4 U724 ( .A(n844), .ZN(n845) );
  INV_X4 U725 ( .A(multinput[20]), .ZN(n844) );
  INV_X4 U726 ( .A(n850), .ZN(n851) );
  INV_X4 U727 ( .A(multinput[23]), .ZN(n850) );
  INV_X4 U728 ( .A(n870), .ZN(n871) );
  INV_X4 U729 ( .A(multinput[33]), .ZN(n870) );
  INV_X4 U730 ( .A(n860), .ZN(n861) );
  INV_X4 U731 ( .A(multinput[28]), .ZN(n860) );
  INV_X4 U732 ( .A(n894), .ZN(n895) );
  INV_X4 U733 ( .A(multinput[45]), .ZN(n894) );
  INV_X4 U734 ( .A(n852), .ZN(n853) );
  INV_X4 U735 ( .A(multinput[24]), .ZN(n852) );
  INV_X4 U736 ( .A(n858), .ZN(n859) );
  INV_X4 U737 ( .A(multinput[27]), .ZN(n858) );
  INV_X4 U738 ( .A(n876), .ZN(n877) );
  INV_X4 U739 ( .A(multinput[36]), .ZN(n876) );
  INV_X4 U740 ( .A(n882), .ZN(n883) );
  INV_X4 U741 ( .A(multinput[39]), .ZN(n882) );
  INV_X4 U742 ( .A(n888), .ZN(n889) );
  INV_X4 U743 ( .A(multinput[42]), .ZN(n888) );
  INV_X4 U744 ( .A(n892), .ZN(n893) );
  INV_X4 U745 ( .A(multinput[44]), .ZN(n892) );
  INV_X4 U746 ( .A(n898), .ZN(n899) );
  INV_X4 U747 ( .A(multinput[47]), .ZN(n898) );
  INV_X4 U748 ( .A(n854), .ZN(n855) );
  INV_X4 U749 ( .A(multinput[25]), .ZN(n854) );
  INV_X4 U750 ( .A(n856), .ZN(n857) );
  INV_X4 U751 ( .A(multinput[26]), .ZN(n856) );
  INV_X4 U752 ( .A(n862), .ZN(n863) );
  INV_X4 U753 ( .A(multinput[29]), .ZN(n862) );
  INV_X4 U754 ( .A(n874), .ZN(n875) );
  INV_X4 U755 ( .A(multinput[35]), .ZN(n874) );
  INV_X4 U756 ( .A(n880), .ZN(n881) );
  INV_X4 U757 ( .A(multinput[38]), .ZN(n880) );
  INV_X4 U758 ( .A(n886), .ZN(n887) );
  INV_X4 U759 ( .A(multinput[41]), .ZN(n886) );
  INV_X4 U760 ( .A(n896), .ZN(n897) );
  INV_X4 U761 ( .A(multinput[46]), .ZN(n896) );
  BUF_X4 U762 ( .A(div_output[0]), .Z(op1[0]) );
  BUF_X4 U763 ( .A(div_output[1]), .Z(op1[1]) );
  BUF_X4 U764 ( .A(div_output[2]), .Z(op1[2]) );
  BUF_X4 U765 ( .A(div_output[3]), .Z(op1[3]) );
  BUF_X4 U766 ( .A(div_output[4]), .Z(op1[4]) );
  BUF_X4 U767 ( .A(div_output[5]), .Z(op1[5]) );
  BUF_X4 U768 ( .A(div_output[6]), .Z(op1[6]) );
  BUF_X4 U769 ( .A(div_output[7]), .Z(op1[7]) );
  BUF_X4 U770 ( .A(div_output[8]), .Z(op1[8]) );
  BUF_X4 U771 ( .A(div_output[9]), .Z(op1[9]) );
  BUF_X4 U772 ( .A(div_output[10]), .Z(op1[10]) );
  BUF_X4 U773 ( .A(div_output[11]), .Z(op1[11]) );
  BUF_X4 U774 ( .A(div_output[12]), .Z(op1[12]) );
  BUF_X4 U775 ( .A(div_output[13]), .Z(op1[13]) );
  BUF_X4 U776 ( .A(div_output[14]), .Z(op1[14]) );
  BUF_X4 U777 ( .A(div_output[15]), .Z(op1[15]) );
  BUF_X4 U778 ( .A(div_output[16]), .Z(op1[16]) );
  BUF_X4 U779 ( .A(div_output[17]), .Z(op1[17]) );
  BUF_X4 U780 ( .A(div_output[18]), .Z(op1[18]) );
  BUF_X4 U781 ( .A(div_output[19]), .Z(op1[19]) );
  BUF_X4 U782 ( .A(div_output[20]), .Z(op1[20]) );
  BUF_X4 U783 ( .A(div_output[21]), .Z(op1[21]) );
  BUF_X4 U784 ( .A(div_output[22]), .Z(op1[22]) );
  BUF_X4 U785 ( .A(div_output[23]), .Z(op1[23]) );
  BUF_X4 U786 ( .A(div_output[24]), .Z(op1[24]) );
  BUF_X4 U787 ( .A(div_output[25]), .Z(op1[25]) );
  BUF_X4 U788 ( .A(div_output[26]), .Z(op1[26]) );
  BUF_X4 U789 ( .A(div_output[27]), .Z(op1[27]) );
  BUF_X4 U790 ( .A(div_output[28]), .Z(op1[28]) );
  BUF_X4 U791 ( .A(div_output[29]), .Z(op1[29]) );
  BUF_X4 U792 ( .A(div_output[30]), .Z(op1[30]) );
  BUF_X4 U793 ( .A(div_output[31]), .Z(op1[31]) );
  BUF_X4 U794 ( .A(div_output[32]), .Z(op1[32]) );
  BUF_X4 U795 ( .A(div_output[33]), .Z(op1[33]) );
  BUF_X4 U796 ( .A(div_output[34]), .Z(op1[34]) );
  BUF_X4 U797 ( .A(div_output[35]), .Z(op1[35]) );
  BUF_X4 U798 ( .A(div_output[36]), .Z(op1[36]) );
  BUF_X4 U799 ( .A(div_output[37]), .Z(op1[37]) );
  BUF_X4 U800 ( .A(div_output[38]), .Z(op1[38]) );
  BUF_X4 U801 ( .A(div_output[39]), .Z(op1[39]) );
  BUF_X4 U802 ( .A(div_output[40]), .Z(op1[40]) );
  BUF_X4 U803 ( .A(div_output[41]), .Z(op1[41]) );
  BUF_X4 U804 ( .A(div_output[42]), .Z(op1[42]) );
  BUF_X4 U805 ( .A(div_output[43]), .Z(op1[43]) );
  BUF_X4 U806 ( .A(div_output[44]), .Z(op1[44]) );
  BUF_X4 U807 ( .A(div_output[45]), .Z(op1[45]) );
  BUF_X4 U808 ( .A(div_output[46]), .Z(op1[46]) );
  BUF_X4 U809 ( .A(div_output[47]), .Z(op1[47]) );
endmodule

